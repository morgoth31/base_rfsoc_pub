----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 05/26/2023 09:36:17 AM
-- Design Name: 
-- Module Name: cos_12table16 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity cos_12table16 is 
    Port ( clk          : in STD_LOGIC;
           angle_12b    : in unsigned (11 downto 0);
           cos_16       : out signed (15 downto 0)
           );
end cos_12table16;


architecture Behavioral of cos_12table16 is
signal angle_12b_conv : std_logic_vector (11 downto 0) ;
begin

angle_12b_conv <= std_logic_vector(angle_12b) ;

process (clk)
begin
    if (rising_edge (clk)) then
        case angle_12b is
        when x"000" => cos_16 <= x"7FFF" ;
        when x"001" => cos_16 <= x"7FFF" ;
        when x"002" => cos_16 <= x"7FFF" ;
        when x"003" => cos_16 <= x"7FFF" ;
        when x"004" => cos_16 <= x"7FFE" ;
        when x"005" => cos_16 <= x"7FFE" ;
        when x"006" => cos_16 <= x"7FFE" ;
        when x"007" => cos_16 <= x"7FFD" ;
        when x"008" => cos_16 <= x"7FFD" ;
        when x"009" => cos_16 <= x"7FFC" ;
        when x"00A" => cos_16 <= x"7FFB" ;
        when x"00B" => cos_16 <= x"7FFA" ;
        when x"00C" => cos_16 <= x"7FF9" ;
        when x"00D" => cos_16 <= x"7FF8" ;
        when x"00E" => cos_16 <= x"7FF7" ;
        when x"00F" => cos_16 <= x"7FF6" ;
        when x"010" => cos_16 <= x"7FF5" ;
        when x"011" => cos_16 <= x"7FF4" ;
        when x"012" => cos_16 <= x"7FF3" ;
        when x"013" => cos_16 <= x"7FF1" ;
        when x"014" => cos_16 <= x"7FF0" ;
        when x"015" => cos_16 <= x"7FEE" ;
        when x"016" => cos_16 <= x"7FEC" ;
        when x"017" => cos_16 <= x"7FEB" ;
        when x"018" => cos_16 <= x"7FE9" ;
        when x"019" => cos_16 <= x"7FE7" ;
        when x"01A" => cos_16 <= x"7FE5" ;
        when x"01B" => cos_16 <= x"7FE3" ;
        when x"01C" => cos_16 <= x"7FE1" ;
        when x"01D" => cos_16 <= x"7FDF" ;
        when x"01E" => cos_16 <= x"7FDC" ;
        when x"01F" => cos_16 <= x"7FDA" ;
        when x"020" => cos_16 <= x"7FD8" ;
        when x"021" => cos_16 <= x"7FD5" ;
        when x"022" => cos_16 <= x"7FD2" ;
        when x"023" => cos_16 <= x"7FD0" ;
        when x"024" => cos_16 <= x"7FCD" ;
        when x"025" => cos_16 <= x"7FCA" ;
        when x"026" => cos_16 <= x"7FC7" ;
        when x"027" => cos_16 <= x"7FC4" ;
        when x"028" => cos_16 <= x"7FC1" ;
        when x"029" => cos_16 <= x"7FBE" ;
        when x"02A" => cos_16 <= x"7FBB" ;
        when x"02B" => cos_16 <= x"7FB8" ;
        when x"02C" => cos_16 <= x"7FB4" ;
        when x"02D" => cos_16 <= x"7FB1" ;
        when x"02E" => cos_16 <= x"7FAD" ;
        when x"02F" => cos_16 <= x"7FAA" ;
        when x"030" => cos_16 <= x"7FA6" ;
        when x"031" => cos_16 <= x"7FA2" ;
        when x"032" => cos_16 <= x"7F9F" ;
        when x"033" => cos_16 <= x"7F9B" ;
        when x"034" => cos_16 <= x"7F97" ;
        when x"035" => cos_16 <= x"7F93" ;
        when x"036" => cos_16 <= x"7F8F" ;
        when x"037" => cos_16 <= x"7F8A" ;
        when x"038" => cos_16 <= x"7F86" ;
        when x"039" => cos_16 <= x"7F82" ;
        when x"03A" => cos_16 <= x"7F7D" ;
        when x"03B" => cos_16 <= x"7F79" ;
        when x"03C" => cos_16 <= x"7F74" ;
        when x"03D" => cos_16 <= x"7F70" ;
        when x"03E" => cos_16 <= x"7F6B" ;
        when x"03F" => cos_16 <= x"7F66" ;
        when x"040" => cos_16 <= x"7F61" ;
        when x"041" => cos_16 <= x"7F5C" ;
        when x"042" => cos_16 <= x"7F57" ;
        when x"043" => cos_16 <= x"7F52" ;
        when x"044" => cos_16 <= x"7F4D" ;
        when x"045" => cos_16 <= x"7F48" ;
        when x"046" => cos_16 <= x"7F42" ;
        when x"047" => cos_16 <= x"7F3D" ;
        when x"048" => cos_16 <= x"7F37" ;
        when x"049" => cos_16 <= x"7F32" ;
        when x"04A" => cos_16 <= x"7F2C" ;
        when x"04B" => cos_16 <= x"7F26" ;
        when x"04C" => cos_16 <= x"7F21" ;
        when x"04D" => cos_16 <= x"7F1B" ;
        when x"04E" => cos_16 <= x"7F15" ;
        when x"04F" => cos_16 <= x"7F0F" ;
        when x"050" => cos_16 <= x"7F09" ;
        when x"051" => cos_16 <= x"7F02" ;
        when x"052" => cos_16 <= x"7EFC" ;
        when x"053" => cos_16 <= x"7EF6" ;
        when x"054" => cos_16 <= x"7EEF" ;
        when x"055" => cos_16 <= x"7EE9" ;
        when x"056" => cos_16 <= x"7EE2" ;
        when x"057" => cos_16 <= x"7EDC" ;
        when x"058" => cos_16 <= x"7ED5" ;
        when x"059" => cos_16 <= x"7ECE" ;
        when x"05A" => cos_16 <= x"7EC7" ;
        when x"05B" => cos_16 <= x"7EC0" ;
        when x"05C" => cos_16 <= x"7EB9" ;
        when x"05D" => cos_16 <= x"7EB2" ;
        when x"05E" => cos_16 <= x"7EAB" ;
        when x"05F" => cos_16 <= x"7EA4" ;
        when x"060" => cos_16 <= x"7E9C" ;
        when x"061" => cos_16 <= x"7E95" ;
        when x"062" => cos_16 <= x"7E8D" ;
        when x"063" => cos_16 <= x"7E86" ;
        when x"064" => cos_16 <= x"7E7E" ;
        when x"065" => cos_16 <= x"7E77" ;
        when x"066" => cos_16 <= x"7E6F" ;
        when x"067" => cos_16 <= x"7E67" ;
        when x"068" => cos_16 <= x"7E5F" ;
        when x"069" => cos_16 <= x"7E57" ;
        when x"06A" => cos_16 <= x"7E4F" ;
        when x"06B" => cos_16 <= x"7E47" ;
        when x"06C" => cos_16 <= x"7E3E" ;
        when x"06D" => cos_16 <= x"7E36" ;
        when x"06E" => cos_16 <= x"7E2E" ;
        when x"06F" => cos_16 <= x"7E25" ;
        when x"070" => cos_16 <= x"7E1D" ;
        when x"071" => cos_16 <= x"7E14" ;
        when x"072" => cos_16 <= x"7E0B" ;
        when x"073" => cos_16 <= x"7E02" ;
        when x"074" => cos_16 <= x"7DFA" ;
        when x"075" => cos_16 <= x"7DF1" ;
        when x"076" => cos_16 <= x"7DE8" ;
        when x"077" => cos_16 <= x"7DDF" ;
        when x"078" => cos_16 <= x"7DD5" ;
        when x"079" => cos_16 <= x"7DCC" ;
        when x"07A" => cos_16 <= x"7DC3" ;
        when x"07B" => cos_16 <= x"7DB9" ;
        when x"07C" => cos_16 <= x"7DB0" ;
        when x"07D" => cos_16 <= x"7DA6" ;
        when x"07E" => cos_16 <= x"7D9D" ;
        when x"07F" => cos_16 <= x"7D93" ;
        when x"080" => cos_16 <= x"7D89" ;
        when x"081" => cos_16 <= x"7D80" ;
        when x"082" => cos_16 <= x"7D76" ;
        when x"083" => cos_16 <= x"7D6C" ;
        when x"084" => cos_16 <= x"7D62" ;
        when x"085" => cos_16 <= x"7D57" ;
        when x"086" => cos_16 <= x"7D4D" ;
        when x"087" => cos_16 <= x"7D43" ;
        when x"088" => cos_16 <= x"7D39" ;
        when x"089" => cos_16 <= x"7D2E" ;
        when x"08A" => cos_16 <= x"7D24" ;
        when x"08B" => cos_16 <= x"7D19" ;
        when x"08C" => cos_16 <= x"7D0E" ;
        when x"08D" => cos_16 <= x"7D04" ;
        when x"08E" => cos_16 <= x"7CF9" ;
        when x"08F" => cos_16 <= x"7CEE" ;
        when x"090" => cos_16 <= x"7CE3" ;
        when x"091" => cos_16 <= x"7CD8" ;
        when x"092" => cos_16 <= x"7CCD" ;
        when x"093" => cos_16 <= x"7CC1" ;
        when x"094" => cos_16 <= x"7CB6" ;
        when x"095" => cos_16 <= x"7CAB" ;
        when x"096" => cos_16 <= x"7C9F" ;
        when x"097" => cos_16 <= x"7C94" ;
        when x"098" => cos_16 <= x"7C88" ;
        when x"099" => cos_16 <= x"7C7D" ;
        when x"09A" => cos_16 <= x"7C71" ;
        when x"09B" => cos_16 <= x"7C65" ;
        when x"09C" => cos_16 <= x"7C59" ;
        when x"09D" => cos_16 <= x"7C4D" ;
        when x"09E" => cos_16 <= x"7C41" ;
        when x"09F" => cos_16 <= x"7C35" ;
        when x"0A0" => cos_16 <= x"7C29" ;
        when x"0A1" => cos_16 <= x"7C1D" ;
        when x"0A2" => cos_16 <= x"7C10" ;
        when x"0A3" => cos_16 <= x"7C04" ;
        when x"0A4" => cos_16 <= x"7BF8" ;
        when x"0A5" => cos_16 <= x"7BEB" ;
        when x"0A6" => cos_16 <= x"7BDE" ;
        when x"0A7" => cos_16 <= x"7BD2" ;
        when x"0A8" => cos_16 <= x"7BC5" ;
        when x"0A9" => cos_16 <= x"7BB8" ;
        when x"0AA" => cos_16 <= x"7BAB" ;
        when x"0AB" => cos_16 <= x"7B9E" ;
        when x"0AC" => cos_16 <= x"7B91" ;
        when x"0AD" => cos_16 <= x"7B84" ;
        when x"0AE" => cos_16 <= x"7B77" ;
        when x"0AF" => cos_16 <= x"7B69" ;
        when x"0B0" => cos_16 <= x"7B5C" ;
        when x"0B1" => cos_16 <= x"7B4F" ;
        when x"0B2" => cos_16 <= x"7B41" ;
        when x"0B3" => cos_16 <= x"7B33" ;
        when x"0B4" => cos_16 <= x"7B26" ;
        when x"0B5" => cos_16 <= x"7B18" ;
        when x"0B6" => cos_16 <= x"7B0A" ;
        when x"0B7" => cos_16 <= x"7AFC" ;
        when x"0B8" => cos_16 <= x"7AEE" ;
        when x"0B9" => cos_16 <= x"7AE0" ;
        when x"0BA" => cos_16 <= x"7AD2" ;
        when x"0BB" => cos_16 <= x"7AC4" ;
        when x"0BC" => cos_16 <= x"7AB6" ;
        when x"0BD" => cos_16 <= x"7AA8" ;
        when x"0BE" => cos_16 <= x"7A99" ;
        when x"0BF" => cos_16 <= x"7A8B" ;
        when x"0C0" => cos_16 <= x"7A7C" ;
        when x"0C1" => cos_16 <= x"7A6D" ;
        when x"0C2" => cos_16 <= x"7A5F" ;
        when x"0C3" => cos_16 <= x"7A50" ;
        when x"0C4" => cos_16 <= x"7A41" ;
        when x"0C5" => cos_16 <= x"7A32" ;
        when x"0C6" => cos_16 <= x"7A23" ;
        when x"0C7" => cos_16 <= x"7A14" ;
        when x"0C8" => cos_16 <= x"7A05" ;
        when x"0C9" => cos_16 <= x"79F6" ;
        when x"0CA" => cos_16 <= x"79E6" ;
        when x"0CB" => cos_16 <= x"79D7" ;
        when x"0CC" => cos_16 <= x"79C8" ;
        when x"0CD" => cos_16 <= x"79B8" ;
        when x"0CE" => cos_16 <= x"79A9" ;
        when x"0CF" => cos_16 <= x"7999" ;
        when x"0D0" => cos_16 <= x"7989" ;
        when x"0D1" => cos_16 <= x"7979" ;
        when x"0D2" => cos_16 <= x"796A" ;
        when x"0D3" => cos_16 <= x"795A" ;
        when x"0D4" => cos_16 <= x"794A" ;
        when x"0D5" => cos_16 <= x"7939" ;
        when x"0D6" => cos_16 <= x"7929" ;
        when x"0D7" => cos_16 <= x"7919" ;
        when x"0D8" => cos_16 <= x"7909" ;
        when x"0D9" => cos_16 <= x"78F8" ;
        when x"0DA" => cos_16 <= x"78E8" ;
        when x"0DB" => cos_16 <= x"78D7" ;
        when x"0DC" => cos_16 <= x"78C7" ;
        when x"0DD" => cos_16 <= x"78B6" ;
        when x"0DE" => cos_16 <= x"78A5" ;
        when x"0DF" => cos_16 <= x"7894" ;
        when x"0E0" => cos_16 <= x"7884" ;
        when x"0E1" => cos_16 <= x"7873" ;
        when x"0E2" => cos_16 <= x"7862" ;
        when x"0E3" => cos_16 <= x"7850" ;
        when x"0E4" => cos_16 <= x"783F" ;
        when x"0E5" => cos_16 <= x"782E" ;
        when x"0E6" => cos_16 <= x"781D" ;
        when x"0E7" => cos_16 <= x"780B" ;
        when x"0E8" => cos_16 <= x"77FA" ;
        when x"0E9" => cos_16 <= x"77E8" ;
        when x"0EA" => cos_16 <= x"77D7" ;
        when x"0EB" => cos_16 <= x"77C5" ;
        when x"0EC" => cos_16 <= x"77B3" ;
        when x"0ED" => cos_16 <= x"77A1" ;
        when x"0EE" => cos_16 <= x"778F" ;
        when x"0EF" => cos_16 <= x"777D" ;
        when x"0F0" => cos_16 <= x"776B" ;
        when x"0F1" => cos_16 <= x"7759" ;
        when x"0F2" => cos_16 <= x"7747" ;
        when x"0F3" => cos_16 <= x"7735" ;
        when x"0F4" => cos_16 <= x"7722" ;
        when x"0F5" => cos_16 <= x"7710" ;
        when x"0F6" => cos_16 <= x"76FE" ;
        when x"0F7" => cos_16 <= x"76EB" ;
        when x"0F8" => cos_16 <= x"76D8" ;
        when x"0F9" => cos_16 <= x"76C6" ;
        when x"0FA" => cos_16 <= x"76B3" ;
        when x"0FB" => cos_16 <= x"76A0" ;
        when x"0FC" => cos_16 <= x"768D" ;
        when x"0FD" => cos_16 <= x"767A" ;
        when x"0FE" => cos_16 <= x"7667" ;
        when x"0FF" => cos_16 <= x"7654" ;
        when x"100" => cos_16 <= x"7641" ;
        when x"101" => cos_16 <= x"762D" ;
        when x"102" => cos_16 <= x"761A" ;
        when x"103" => cos_16 <= x"7607" ;
        when x"104" => cos_16 <= x"75F3" ;
        when x"105" => cos_16 <= x"75E0" ;
        when x"106" => cos_16 <= x"75CC" ;
        when x"107" => cos_16 <= x"75B8" ;
        when x"108" => cos_16 <= x"75A5" ;
        when x"109" => cos_16 <= x"7591" ;
        when x"10A" => cos_16 <= x"757D" ;
        when x"10B" => cos_16 <= x"7569" ;
        when x"10C" => cos_16 <= x"7555" ;
        when x"10D" => cos_16 <= x"7541" ;
        when x"10E" => cos_16 <= x"752D" ;
        when x"10F" => cos_16 <= x"7518" ;
        when x"110" => cos_16 <= x"7504" ;
        when x"111" => cos_16 <= x"74F0" ;
        when x"112" => cos_16 <= x"74DB" ;
        when x"113" => cos_16 <= x"74C6" ;
        when x"114" => cos_16 <= x"74B2" ;
        when x"115" => cos_16 <= x"749D" ;
        when x"116" => cos_16 <= x"7488" ;
        when x"117" => cos_16 <= x"7474" ;
        when x"118" => cos_16 <= x"745F" ;
        when x"119" => cos_16 <= x"744A" ;
        when x"11A" => cos_16 <= x"7435" ;
        when x"11B" => cos_16 <= x"7420" ;
        when x"11C" => cos_16 <= x"740A" ;
        when x"11D" => cos_16 <= x"73F5" ;
        when x"11E" => cos_16 <= x"73E0" ;
        when x"11F" => cos_16 <= x"73CA" ;
        when x"120" => cos_16 <= x"73B5" ;
        when x"121" => cos_16 <= x"739F" ;
        when x"122" => cos_16 <= x"738A" ;
        when x"123" => cos_16 <= x"7374" ;
        when x"124" => cos_16 <= x"735E" ;
        when x"125" => cos_16 <= x"7349" ;
        when x"126" => cos_16 <= x"7333" ;
        when x"127" => cos_16 <= x"731D" ;
        when x"128" => cos_16 <= x"7307" ;
        when x"129" => cos_16 <= x"72F1" ;
        when x"12A" => cos_16 <= x"72DB" ;
        when x"12B" => cos_16 <= x"72C4" ;
        when x"12C" => cos_16 <= x"72AE" ;
        when x"12D" => cos_16 <= x"7298" ;
        when x"12E" => cos_16 <= x"7281" ;
        when x"12F" => cos_16 <= x"726B" ;
        when x"130" => cos_16 <= x"7254" ;
        when x"131" => cos_16 <= x"723E" ;
        when x"132" => cos_16 <= x"7227" ;
        when x"133" => cos_16 <= x"7210" ;
        when x"134" => cos_16 <= x"71F9" ;
        when x"135" => cos_16 <= x"71E2" ;
        when x"136" => cos_16 <= x"71CB" ;
        when x"137" => cos_16 <= x"71B4" ;
        when x"138" => cos_16 <= x"719D" ;
        when x"139" => cos_16 <= x"7186" ;
        when x"13A" => cos_16 <= x"716F" ;
        when x"13B" => cos_16 <= x"7158" ;
        when x"13C" => cos_16 <= x"7140" ;
        when x"13D" => cos_16 <= x"7129" ;
        when x"13E" => cos_16 <= x"7111" ;
        when x"13F" => cos_16 <= x"70FA" ;
        when x"140" => cos_16 <= x"70E2" ;
        when x"141" => cos_16 <= x"70CA" ;
        when x"142" => cos_16 <= x"70B2" ;
        when x"143" => cos_16 <= x"709B" ;
        when x"144" => cos_16 <= x"7083" ;
        when x"145" => cos_16 <= x"706B" ;
        when x"146" => cos_16 <= x"7053" ;
        when x"147" => cos_16 <= x"703A" ;
        when x"148" => cos_16 <= x"7022" ;
        when x"149" => cos_16 <= x"700A" ;
        when x"14A" => cos_16 <= x"6FF2" ;
        when x"14B" => cos_16 <= x"6FD9" ;
        when x"14C" => cos_16 <= x"6FC1" ;
        when x"14D" => cos_16 <= x"6FA8" ;
        when x"14E" => cos_16 <= x"6F90" ;
        when x"14F" => cos_16 <= x"6F77" ;
        when x"150" => cos_16 <= x"6F5E" ;
        when x"151" => cos_16 <= x"6F45" ;
        when x"152" => cos_16 <= x"6F2C" ;
        when x"153" => cos_16 <= x"6F14" ;
        when x"154" => cos_16 <= x"6EFB" ;
        when x"155" => cos_16 <= x"6EE1" ;
        when x"156" => cos_16 <= x"6EC8" ;
        when x"157" => cos_16 <= x"6EAF" ;
        when x"158" => cos_16 <= x"6E96" ;
        when x"159" => cos_16 <= x"6E7C" ;
        when x"15A" => cos_16 <= x"6E63" ;
        when x"15B" => cos_16 <= x"6E4A" ;
        when x"15C" => cos_16 <= x"6E30" ;
        when x"15D" => cos_16 <= x"6E16" ;
        when x"15E" => cos_16 <= x"6DFD" ;
        when x"15F" => cos_16 <= x"6DE3" ;
        when x"160" => cos_16 <= x"6DC9" ;
        when x"161" => cos_16 <= x"6DAF" ;
        when x"162" => cos_16 <= x"6D95" ;
        when x"163" => cos_16 <= x"6D7B" ;
        when x"164" => cos_16 <= x"6D61" ;
        when x"165" => cos_16 <= x"6D47" ;
        when x"166" => cos_16 <= x"6D2D" ;
        when x"167" => cos_16 <= x"6D13" ;
        when x"168" => cos_16 <= x"6CF8" ;
        when x"169" => cos_16 <= x"6CDE" ;
        when x"16A" => cos_16 <= x"6CC3" ;
        when x"16B" => cos_16 <= x"6CA9" ;
        when x"16C" => cos_16 <= x"6C8E" ;
        when x"16D" => cos_16 <= x"6C74" ;
        when x"16E" => cos_16 <= x"6C59" ;
        when x"16F" => cos_16 <= x"6C3E" ;
        when x"170" => cos_16 <= x"6C23" ;
        when x"171" => cos_16 <= x"6C08" ;
        when x"172" => cos_16 <= x"6BED" ;
        when x"173" => cos_16 <= x"6BD2" ;
        when x"174" => cos_16 <= x"6BB7" ;
        when x"175" => cos_16 <= x"6B9C" ;
        when x"176" => cos_16 <= x"6B81" ;
        when x"177" => cos_16 <= x"6B65" ;
        when x"178" => cos_16 <= x"6B4A" ;
        when x"179" => cos_16 <= x"6B2F" ;
        when x"17A" => cos_16 <= x"6B13" ;
        when x"17B" => cos_16 <= x"6AF8" ;
        when x"17C" => cos_16 <= x"6ADC" ;
        when x"17D" => cos_16 <= x"6AC0" ;
        when x"17E" => cos_16 <= x"6AA4" ;
        when x"17F" => cos_16 <= x"6A89" ;
        when x"180" => cos_16 <= x"6A6D" ;
        when x"181" => cos_16 <= x"6A51" ;
        when x"182" => cos_16 <= x"6A35" ;
        when x"183" => cos_16 <= x"6A19" ;
        when x"184" => cos_16 <= x"69FD" ;
        when x"185" => cos_16 <= x"69E0" ;
        when x"186" => cos_16 <= x"69C4" ;
        when x"187" => cos_16 <= x"69A8" ;
        when x"188" => cos_16 <= x"698B" ;
        when x"189" => cos_16 <= x"696F" ;
        when x"18A" => cos_16 <= x"6952" ;
        when x"18B" => cos_16 <= x"6936" ;
        when x"18C" => cos_16 <= x"6919" ;
        when x"18D" => cos_16 <= x"68FC" ;
        when x"18E" => cos_16 <= x"68E0" ;
        when x"18F" => cos_16 <= x"68C3" ;
        when x"190" => cos_16 <= x"68A6" ;
        when x"191" => cos_16 <= x"6889" ;
        when x"192" => cos_16 <= x"686C" ;
        when x"193" => cos_16 <= x"684F" ;
        when x"194" => cos_16 <= x"6832" ;
        when x"195" => cos_16 <= x"6814" ;
        when x"196" => cos_16 <= x"67F7" ;
        when x"197" => cos_16 <= x"67DA" ;
        when x"198" => cos_16 <= x"67BC" ;
        when x"199" => cos_16 <= x"679F" ;
        when x"19A" => cos_16 <= x"6781" ;
        when x"19B" => cos_16 <= x"6764" ;
        when x"19C" => cos_16 <= x"6746" ;
        when x"19D" => cos_16 <= x"6728" ;
        when x"19E" => cos_16 <= x"670A" ;
        when x"19F" => cos_16 <= x"66ED" ;
        when x"1A0" => cos_16 <= x"66CF" ;
        when x"1A1" => cos_16 <= x"66B1" ;
        when x"1A2" => cos_16 <= x"6693" ;
        when x"1A3" => cos_16 <= x"6675" ;
        when x"1A4" => cos_16 <= x"6656" ;
        when x"1A5" => cos_16 <= x"6638" ;
        when x"1A6" => cos_16 <= x"661A" ;
        when x"1A7" => cos_16 <= x"65FC" ;
        when x"1A8" => cos_16 <= x"65DD" ;
        when x"1A9" => cos_16 <= x"65BF" ;
        when x"1AA" => cos_16 <= x"65A0" ;
        when x"1AB" => cos_16 <= x"6582" ;
        when x"1AC" => cos_16 <= x"6563" ;
        when x"1AD" => cos_16 <= x"6544" ;
        when x"1AE" => cos_16 <= x"6525" ;
        when x"1AF" => cos_16 <= x"6507" ;
        when x"1B0" => cos_16 <= x"64E8" ;
        when x"1B1" => cos_16 <= x"64C9" ;
        when x"1B2" => cos_16 <= x"64AA" ;
        when x"1B3" => cos_16 <= x"648B" ;
        when x"1B4" => cos_16 <= x"646C" ;
        when x"1B5" => cos_16 <= x"644C" ;
        when x"1B6" => cos_16 <= x"642D" ;
        when x"1B7" => cos_16 <= x"640E" ;
        when x"1B8" => cos_16 <= x"63EE" ;
        when x"1B9" => cos_16 <= x"63CF" ;
        when x"1BA" => cos_16 <= x"63AF" ;
        when x"1BB" => cos_16 <= x"6390" ;
        when x"1BC" => cos_16 <= x"6370" ;
        when x"1BD" => cos_16 <= x"6351" ;
        when x"1BE" => cos_16 <= x"6331" ;
        when x"1BF" => cos_16 <= x"6311" ;
        when x"1C0" => cos_16 <= x"62F1" ;
        when x"1C1" => cos_16 <= x"62D1" ;
        when x"1C2" => cos_16 <= x"62B1" ;
        when x"1C3" => cos_16 <= x"6291" ;
        when x"1C4" => cos_16 <= x"6271" ;
        when x"1C5" => cos_16 <= x"6251" ;
        when x"1C6" => cos_16 <= x"6231" ;
        when x"1C7" => cos_16 <= x"6211" ;
        when x"1C8" => cos_16 <= x"61F0" ;
        when x"1C9" => cos_16 <= x"61D0" ;
        when x"1CA" => cos_16 <= x"61AF" ;
        when x"1CB" => cos_16 <= x"618F" ;
        when x"1CC" => cos_16 <= x"616E" ;
        when x"1CD" => cos_16 <= x"614E" ;
        when x"1CE" => cos_16 <= x"612D" ;
        when x"1CF" => cos_16 <= x"610C" ;
        when x"1D0" => cos_16 <= x"60EB" ;
        when x"1D1" => cos_16 <= x"60CB" ;
        when x"1D2" => cos_16 <= x"60AA" ;
        when x"1D3" => cos_16 <= x"6089" ;
        when x"1D4" => cos_16 <= x"6068" ;
        when x"1D5" => cos_16 <= x"6047" ;
        when x"1D6" => cos_16 <= x"6025" ;
        when x"1D7" => cos_16 <= x"6004" ;
        when x"1D8" => cos_16 <= x"5FE3" ;
        when x"1D9" => cos_16 <= x"5FC2" ;
        when x"1DA" => cos_16 <= x"5FA0" ;
        when x"1DB" => cos_16 <= x"5F7F" ;
        when x"1DC" => cos_16 <= x"5F5D" ;
        when x"1DD" => cos_16 <= x"5F3C" ;
        when x"1DE" => cos_16 <= x"5F1A" ;
        when x"1DF" => cos_16 <= x"5EF8" ;
        when x"1E0" => cos_16 <= x"5ED7" ;
        when x"1E1" => cos_16 <= x"5EB5" ;
        when x"1E2" => cos_16 <= x"5E93" ;
        when x"1E3" => cos_16 <= x"5E71" ;
        when x"1E4" => cos_16 <= x"5E4F" ;
        when x"1E5" => cos_16 <= x"5E2D" ;
        when x"1E6" => cos_16 <= x"5E0B" ;
        when x"1E7" => cos_16 <= x"5DE9" ;
        when x"1E8" => cos_16 <= x"5DC7" ;
        when x"1E9" => cos_16 <= x"5DA5" ;
        when x"1EA" => cos_16 <= x"5D82" ;
        when x"1EB" => cos_16 <= x"5D60" ;
        when x"1EC" => cos_16 <= x"5D3E" ;
        when x"1ED" => cos_16 <= x"5D1B" ;
        when x"1EE" => cos_16 <= x"5CF9" ;
        when x"1EF" => cos_16 <= x"5CD6" ;
        when x"1F0" => cos_16 <= x"5CB3" ;
        when x"1F1" => cos_16 <= x"5C91" ;
        when x"1F2" => cos_16 <= x"5C6E" ;
        when x"1F3" => cos_16 <= x"5C4B" ;
        when x"1F4" => cos_16 <= x"5C28" ;
        when x"1F5" => cos_16 <= x"5C05" ;
        when x"1F6" => cos_16 <= x"5BE2" ;
        when x"1F7" => cos_16 <= x"5BBF" ;
        when x"1F8" => cos_16 <= x"5B9C" ;
        when x"1F9" => cos_16 <= x"5B79" ;
        when x"1FA" => cos_16 <= x"5B56" ;
        when x"1FB" => cos_16 <= x"5B33" ;
        when x"1FC" => cos_16 <= x"5B0F" ;
        when x"1FD" => cos_16 <= x"5AEC" ;
        when x"1FE" => cos_16 <= x"5AC9" ;
        when x"1FF" => cos_16 <= x"5AA5" ;
        when x"200" => cos_16 <= x"5A82" ;
        when x"201" => cos_16 <= x"5A5E" ;
        when x"202" => cos_16 <= x"5A3B" ;
        when x"203" => cos_16 <= x"5A17" ;
        when x"204" => cos_16 <= x"59F3" ;
        when x"205" => cos_16 <= x"59CF" ;
        when x"206" => cos_16 <= x"59AC" ;
        when x"207" => cos_16 <= x"5988" ;
        when x"208" => cos_16 <= x"5964" ;
        when x"209" => cos_16 <= x"5940" ;
        when x"20A" => cos_16 <= x"591C" ;
        when x"20B" => cos_16 <= x"58F8" ;
        when x"20C" => cos_16 <= x"58D3" ;
        when x"20D" => cos_16 <= x"58AF" ;
        when x"20E" => cos_16 <= x"588B" ;
        when x"20F" => cos_16 <= x"5867" ;
        when x"210" => cos_16 <= x"5842" ;
        when x"211" => cos_16 <= x"581E" ;
        when x"212" => cos_16 <= x"57F9" ;
        when x"213" => cos_16 <= x"57D5" ;
        when x"214" => cos_16 <= x"57B0" ;
        when x"215" => cos_16 <= x"578B" ;
        when x"216" => cos_16 <= x"5767" ;
        when x"217" => cos_16 <= x"5742" ;
        when x"218" => cos_16 <= x"571D" ;
        when x"219" => cos_16 <= x"56F8" ;
        when x"21A" => cos_16 <= x"56D3" ;
        when x"21B" => cos_16 <= x"56AF" ;
        when x"21C" => cos_16 <= x"568A" ;
        when x"21D" => cos_16 <= x"5664" ;
        when x"21E" => cos_16 <= x"563F" ;
        when x"21F" => cos_16 <= x"561A" ;
        when x"220" => cos_16 <= x"55F5" ;
        when x"221" => cos_16 <= x"55D0" ;
        when x"222" => cos_16 <= x"55AA" ;
        when x"223" => cos_16 <= x"5585" ;
        when x"224" => cos_16 <= x"5560" ;
        when x"225" => cos_16 <= x"553A" ;
        when x"226" => cos_16 <= x"5515" ;
        when x"227" => cos_16 <= x"54EF" ;
        when x"228" => cos_16 <= x"54C9" ;
        when x"229" => cos_16 <= x"54A4" ;
        when x"22A" => cos_16 <= x"547E" ;
        when x"22B" => cos_16 <= x"5458" ;
        when x"22C" => cos_16 <= x"5432" ;
        when x"22D" => cos_16 <= x"540C" ;
        when x"22E" => cos_16 <= x"53E7" ;
        when x"22F" => cos_16 <= x"53C1" ;
        when x"230" => cos_16 <= x"539B" ;
        when x"231" => cos_16 <= x"5374" ;
        when x"232" => cos_16 <= x"534E" ;
        when x"233" => cos_16 <= x"5328" ;
        when x"234" => cos_16 <= x"5302" ;
        when x"235" => cos_16 <= x"52DC" ;
        when x"236" => cos_16 <= x"52B5" ;
        when x"237" => cos_16 <= x"528F" ;
        when x"238" => cos_16 <= x"5268" ;
        when x"239" => cos_16 <= x"5242" ;
        when x"23A" => cos_16 <= x"521B" ;
        when x"23B" => cos_16 <= x"51F5" ;
        when x"23C" => cos_16 <= x"51CE" ;
        when x"23D" => cos_16 <= x"51A8" ;
        when x"23E" => cos_16 <= x"5181" ;
        when x"23F" => cos_16 <= x"515A" ;
        when x"240" => cos_16 <= x"5133" ;
        when x"241" => cos_16 <= x"510C" ;
        when x"242" => cos_16 <= x"50E5" ;
        when x"243" => cos_16 <= x"50BE" ;
        when x"244" => cos_16 <= x"5097" ;
        when x"245" => cos_16 <= x"5070" ;
        when x"246" => cos_16 <= x"5049" ;
        when x"247" => cos_16 <= x"5022" ;
        when x"248" => cos_16 <= x"4FFB" ;
        when x"249" => cos_16 <= x"4FD4" ;
        when x"24A" => cos_16 <= x"4FAC" ;
        when x"24B" => cos_16 <= x"4F85" ;
        when x"24C" => cos_16 <= x"4F5D" ;
        when x"24D" => cos_16 <= x"4F36" ;
        when x"24E" => cos_16 <= x"4F0E" ;
        when x"24F" => cos_16 <= x"4EE7" ;
        when x"250" => cos_16 <= x"4EBF" ;
        when x"251" => cos_16 <= x"4E98" ;
        when x"252" => cos_16 <= x"4E70" ;
        when x"253" => cos_16 <= x"4E48" ;
        when x"254" => cos_16 <= x"4E20" ;
        when x"255" => cos_16 <= x"4DF9" ;
        when x"256" => cos_16 <= x"4DD1" ;
        when x"257" => cos_16 <= x"4DA9" ;
        when x"258" => cos_16 <= x"4D81" ;
        when x"259" => cos_16 <= x"4D59" ;
        when x"25A" => cos_16 <= x"4D31" ;
        when x"25B" => cos_16 <= x"4D09" ;
        when x"25C" => cos_16 <= x"4CE0" ;
        when x"25D" => cos_16 <= x"4CB8" ;
        when x"25E" => cos_16 <= x"4C90" ;
        when x"25F" => cos_16 <= x"4C68" ;
        when x"260" => cos_16 <= x"4C3F" ;
        when x"261" => cos_16 <= x"4C17" ;
        when x"262" => cos_16 <= x"4BEE" ;
        when x"263" => cos_16 <= x"4BC6" ;
        when x"264" => cos_16 <= x"4B9D" ;
        when x"265" => cos_16 <= x"4B75" ;
        when x"266" => cos_16 <= x"4B4C" ;
        when x"267" => cos_16 <= x"4B24" ;
        when x"268" => cos_16 <= x"4AFB" ;
        when x"269" => cos_16 <= x"4AD2" ;
        when x"26A" => cos_16 <= x"4AA9" ;
        when x"26B" => cos_16 <= x"4A80" ;
        when x"26C" => cos_16 <= x"4A58" ;
        when x"26D" => cos_16 <= x"4A2F" ;
        when x"26E" => cos_16 <= x"4A06" ;
        when x"26F" => cos_16 <= x"49DD" ;
        when x"270" => cos_16 <= x"49B4" ;
        when x"271" => cos_16 <= x"498A" ;
        when x"272" => cos_16 <= x"4961" ;
        when x"273" => cos_16 <= x"4938" ;
        when x"274" => cos_16 <= x"490F" ;
        when x"275" => cos_16 <= x"48E5" ;
        when x"276" => cos_16 <= x"48BC" ;
        when x"277" => cos_16 <= x"4893" ;
        when x"278" => cos_16 <= x"4869" ;
        when x"279" => cos_16 <= x"4840" ;
        when x"27A" => cos_16 <= x"4816" ;
        when x"27B" => cos_16 <= x"47ED" ;
        when x"27C" => cos_16 <= x"47C3" ;
        when x"27D" => cos_16 <= x"479A" ;
        when x"27E" => cos_16 <= x"4770" ;
        when x"27F" => cos_16 <= x"4746" ;
        when x"280" => cos_16 <= x"471C" ;
        when x"281" => cos_16 <= x"46F3" ;
        when x"282" => cos_16 <= x"46C9" ;
        when x"283" => cos_16 <= x"469F" ;
        when x"284" => cos_16 <= x"4675" ;
        when x"285" => cos_16 <= x"464B" ;
        when x"286" => cos_16 <= x"4621" ;
        when x"287" => cos_16 <= x"45F7" ;
        when x"288" => cos_16 <= x"45CD" ;
        when x"289" => cos_16 <= x"45A3" ;
        when x"28A" => cos_16 <= x"4578" ;
        when x"28B" => cos_16 <= x"454E" ;
        when x"28C" => cos_16 <= x"4524" ;
        when x"28D" => cos_16 <= x"44F9" ;
        when x"28E" => cos_16 <= x"44CF" ;
        when x"28F" => cos_16 <= x"44A5" ;
        when x"290" => cos_16 <= x"447A" ;
        when x"291" => cos_16 <= x"4450" ;
        when x"292" => cos_16 <= x"4425" ;
        when x"293" => cos_16 <= x"43FB" ;
        when x"294" => cos_16 <= x"43D0" ;
        when x"295" => cos_16 <= x"43A5" ;
        when x"296" => cos_16 <= x"437B" ;
        when x"297" => cos_16 <= x"4350" ;
        when x"298" => cos_16 <= x"4325" ;
        when x"299" => cos_16 <= x"42FA" ;
        when x"29A" => cos_16 <= x"42D0" ;
        when x"29B" => cos_16 <= x"42A5" ;
        when x"29C" => cos_16 <= x"427A" ;
        when x"29D" => cos_16 <= x"424F" ;
        when x"29E" => cos_16 <= x"4224" ;
        when x"29F" => cos_16 <= x"41F9" ;
        when x"2A0" => cos_16 <= x"41CE" ;
        when x"2A1" => cos_16 <= x"41A2" ;
        when x"2A2" => cos_16 <= x"4177" ;
        when x"2A3" => cos_16 <= x"414C" ;
        when x"2A4" => cos_16 <= x"4121" ;
        when x"2A5" => cos_16 <= x"40F6" ;
        when x"2A6" => cos_16 <= x"40CA" ;
        when x"2A7" => cos_16 <= x"409F" ;
        when x"2A8" => cos_16 <= x"4073" ;
        when x"2A9" => cos_16 <= x"4048" ;
        when x"2AA" => cos_16 <= x"401D" ;
        when x"2AB" => cos_16 <= x"3FF1" ;
        when x"2AC" => cos_16 <= x"3FC5" ;
        when x"2AD" => cos_16 <= x"3F9A" ;
        when x"2AE" => cos_16 <= x"3F6E" ;
        when x"2AF" => cos_16 <= x"3F43" ;
        when x"2B0" => cos_16 <= x"3F17" ;
        when x"2B1" => cos_16 <= x"3EEB" ;
        when x"2B2" => cos_16 <= x"3EBF" ;
        when x"2B3" => cos_16 <= x"3E93" ;
        when x"2B4" => cos_16 <= x"3E68" ;
        when x"2B5" => cos_16 <= x"3E3C" ;
        when x"2B6" => cos_16 <= x"3E10" ;
        when x"2B7" => cos_16 <= x"3DE4" ;
        when x"2B8" => cos_16 <= x"3DB8" ;
        when x"2B9" => cos_16 <= x"3D8C" ;
        when x"2BA" => cos_16 <= x"3D60" ;
        when x"2BB" => cos_16 <= x"3D33" ;
        when x"2BC" => cos_16 <= x"3D07" ;
        when x"2BD" => cos_16 <= x"3CDB" ;
        when x"2BE" => cos_16 <= x"3CAF" ;
        when x"2BF" => cos_16 <= x"3C83" ;
        when x"2C0" => cos_16 <= x"3C56" ;
        when x"2C1" => cos_16 <= x"3C2A" ;
        when x"2C2" => cos_16 <= x"3BFE" ;
        when x"2C3" => cos_16 <= x"3BD1" ;
        when x"2C4" => cos_16 <= x"3BA5" ;
        when x"2C5" => cos_16 <= x"3B78" ;
        when x"2C6" => cos_16 <= x"3B4C" ;
        when x"2C7" => cos_16 <= x"3B1F" ;
        when x"2C8" => cos_16 <= x"3AF2" ;
        when x"2C9" => cos_16 <= x"3AC6" ;
        when x"2CA" => cos_16 <= x"3A99" ;
        when x"2CB" => cos_16 <= x"3A6C" ;
        when x"2CC" => cos_16 <= x"3A40" ;
        when x"2CD" => cos_16 <= x"3A13" ;
        when x"2CE" => cos_16 <= x"39E6" ;
        when x"2CF" => cos_16 <= x"39B9" ;
        when x"2D0" => cos_16 <= x"398C" ;
        when x"2D1" => cos_16 <= x"3960" ;
        when x"2D2" => cos_16 <= x"3933" ;
        when x"2D3" => cos_16 <= x"3906" ;
        when x"2D4" => cos_16 <= x"38D9" ;
        when x"2D5" => cos_16 <= x"38AB" ;
        when x"2D6" => cos_16 <= x"387E" ;
        when x"2D7" => cos_16 <= x"3851" ;
        when x"2D8" => cos_16 <= x"3824" ;
        when x"2D9" => cos_16 <= x"37F7" ;
        when x"2DA" => cos_16 <= x"37CA" ;
        when x"2DB" => cos_16 <= x"379C" ;
        when x"2DC" => cos_16 <= x"376F" ;
        when x"2DD" => cos_16 <= x"3742" ;
        when x"2DE" => cos_16 <= x"3715" ;
        when x"2DF" => cos_16 <= x"36E7" ;
        when x"2E0" => cos_16 <= x"36BA" ;
        when x"2E1" => cos_16 <= x"368C" ;
        when x"2E2" => cos_16 <= x"365F" ;
        when x"2E3" => cos_16 <= x"3631" ;
        when x"2E4" => cos_16 <= x"3604" ;
        when x"2E5" => cos_16 <= x"35D6" ;
        when x"2E6" => cos_16 <= x"35A8" ;
        when x"2E7" => cos_16 <= x"357B" ;
        when x"2E8" => cos_16 <= x"354D" ;
        when x"2E9" => cos_16 <= x"351F" ;
        when x"2EA" => cos_16 <= x"34F2" ;
        when x"2EB" => cos_16 <= x"34C4" ;
        when x"2EC" => cos_16 <= x"3496" ;
        when x"2ED" => cos_16 <= x"3468" ;
        when x"2EE" => cos_16 <= x"343A" ;
        when x"2EF" => cos_16 <= x"340C" ;
        when x"2F0" => cos_16 <= x"33DF" ;
        when x"2F1" => cos_16 <= x"33B1" ;
        when x"2F2" => cos_16 <= x"3383" ;
        when x"2F3" => cos_16 <= x"3355" ;
        when x"2F4" => cos_16 <= x"3326" ;
        when x"2F5" => cos_16 <= x"32F8" ;
        when x"2F6" => cos_16 <= x"32CA" ;
        when x"2F7" => cos_16 <= x"329C" ;
        when x"2F8" => cos_16 <= x"326E" ;
        when x"2F9" => cos_16 <= x"3240" ;
        when x"2FA" => cos_16 <= x"3211" ;
        when x"2FB" => cos_16 <= x"31E3" ;
        when x"2FC" => cos_16 <= x"31B5" ;
        when x"2FD" => cos_16 <= x"3187" ;
        when x"2FE" => cos_16 <= x"3158" ;
        when x"2FF" => cos_16 <= x"312A" ;
        when x"300" => cos_16 <= x"30FB" ;
        when x"301" => cos_16 <= x"30CD" ;
        when x"302" => cos_16 <= x"309E" ;
        when x"303" => cos_16 <= x"3070" ;
        when x"304" => cos_16 <= x"3041" ;
        when x"305" => cos_16 <= x"3013" ;
        when x"306" => cos_16 <= x"2FE4" ;
        when x"307" => cos_16 <= x"2FB6" ;
        when x"308" => cos_16 <= x"2F87" ;
        when x"309" => cos_16 <= x"2F58" ;
        when x"30A" => cos_16 <= x"2F2A" ;
        when x"30B" => cos_16 <= x"2EFB" ;
        when x"30C" => cos_16 <= x"2ECC" ;
        when x"30D" => cos_16 <= x"2E9D" ;
        when x"30E" => cos_16 <= x"2E6E" ;
        when x"30F" => cos_16 <= x"2E40" ;
        when x"310" => cos_16 <= x"2E11" ;
        when x"311" => cos_16 <= x"2DE2" ;
        when x"312" => cos_16 <= x"2DB3" ;
        when x"313" => cos_16 <= x"2D84" ;
        when x"314" => cos_16 <= x"2D55" ;
        when x"315" => cos_16 <= x"2D26" ;
        when x"316" => cos_16 <= x"2CF7" ;
        when x"317" => cos_16 <= x"2CC8" ;
        when x"318" => cos_16 <= x"2C99" ;
        when x"319" => cos_16 <= x"2C6A" ;
        when x"31A" => cos_16 <= x"2C3A" ;
        when x"31B" => cos_16 <= x"2C0B" ;
        when x"31C" => cos_16 <= x"2BDC" ;
        when x"31D" => cos_16 <= x"2BAD" ;
        when x"31E" => cos_16 <= x"2B7D" ;
        when x"31F" => cos_16 <= x"2B4E" ;
        when x"320" => cos_16 <= x"2B1F" ;
        when x"321" => cos_16 <= x"2AF0" ;
        when x"322" => cos_16 <= x"2AC0" ;
        when x"323" => cos_16 <= x"2A91" ;
        when x"324" => cos_16 <= x"2A61" ;
        when x"325" => cos_16 <= x"2A32" ;
        when x"326" => cos_16 <= x"2A02" ;
        when x"327" => cos_16 <= x"29D3" ;
        when x"328" => cos_16 <= x"29A3" ;
        when x"329" => cos_16 <= x"2974" ;
        when x"32A" => cos_16 <= x"2944" ;
        when x"32B" => cos_16 <= x"2915" ;
        when x"32C" => cos_16 <= x"28E5" ;
        when x"32D" => cos_16 <= x"28B5" ;
        when x"32E" => cos_16 <= x"2886" ;
        when x"32F" => cos_16 <= x"2856" ;
        when x"330" => cos_16 <= x"2826" ;
        when x"331" => cos_16 <= x"27F7" ;
        when x"332" => cos_16 <= x"27C7" ;
        when x"333" => cos_16 <= x"2797" ;
        when x"334" => cos_16 <= x"2767" ;
        when x"335" => cos_16 <= x"2737" ;
        when x"336" => cos_16 <= x"2708" ;
        when x"337" => cos_16 <= x"26D8" ;
        when x"338" => cos_16 <= x"26A8" ;
        when x"339" => cos_16 <= x"2678" ;
        when x"33A" => cos_16 <= x"2648" ;
        when x"33B" => cos_16 <= x"2618" ;
        when x"33C" => cos_16 <= x"25E8" ;
        when x"33D" => cos_16 <= x"25B8" ;
        when x"33E" => cos_16 <= x"2588" ;
        when x"33F" => cos_16 <= x"2558" ;
        when x"340" => cos_16 <= x"2528" ;
        when x"341" => cos_16 <= x"24F8" ;
        when x"342" => cos_16 <= x"24C8" ;
        when x"343" => cos_16 <= x"2497" ;
        when x"344" => cos_16 <= x"2467" ;
        when x"345" => cos_16 <= x"2437" ;
        when x"346" => cos_16 <= x"2407" ;
        when x"347" => cos_16 <= x"23D7" ;
        when x"348" => cos_16 <= x"23A6" ;
        when x"349" => cos_16 <= x"2376" ;
        when x"34A" => cos_16 <= x"2346" ;
        when x"34B" => cos_16 <= x"2315" ;
        when x"34C" => cos_16 <= x"22E5" ;
        when x"34D" => cos_16 <= x"22B5" ;
        when x"34E" => cos_16 <= x"2284" ;
        when x"34F" => cos_16 <= x"2254" ;
        when x"350" => cos_16 <= x"2223" ;
        when x"351" => cos_16 <= x"21F3" ;
        when x"352" => cos_16 <= x"21C2" ;
        when x"353" => cos_16 <= x"2192" ;
        when x"354" => cos_16 <= x"2161" ;
        when x"355" => cos_16 <= x"2131" ;
        when x"356" => cos_16 <= x"2100" ;
        when x"357" => cos_16 <= x"20D0" ;
        when x"358" => cos_16 <= x"209F" ;
        when x"359" => cos_16 <= x"206F" ;
        when x"35A" => cos_16 <= x"203E" ;
        when x"35B" => cos_16 <= x"200D" ;
        when x"35C" => cos_16 <= x"1FDD" ;
        when x"35D" => cos_16 <= x"1FAC" ;
        when x"35E" => cos_16 <= x"1F7B" ;
        when x"35F" => cos_16 <= x"1F4A" ;
        when x"360" => cos_16 <= x"1F1A" ;
        when x"361" => cos_16 <= x"1EE9" ;
        when x"362" => cos_16 <= x"1EB8" ;
        when x"363" => cos_16 <= x"1E87" ;
        when x"364" => cos_16 <= x"1E57" ;
        when x"365" => cos_16 <= x"1E26" ;
        when x"366" => cos_16 <= x"1DF5" ;
        when x"367" => cos_16 <= x"1DC4" ;
        when x"368" => cos_16 <= x"1D93" ;
        when x"369" => cos_16 <= x"1D62" ;
        when x"36A" => cos_16 <= x"1D31" ;
        when x"36B" => cos_16 <= x"1D00" ;
        when x"36C" => cos_16 <= x"1CCF" ;
        when x"36D" => cos_16 <= x"1C9E" ;
        when x"36E" => cos_16 <= x"1C6D" ;
        when x"36F" => cos_16 <= x"1C3C" ;
        when x"370" => cos_16 <= x"1C0B" ;
        when x"371" => cos_16 <= x"1BDA" ;
        when x"372" => cos_16 <= x"1BA9" ;
        when x"373" => cos_16 <= x"1B78" ;
        when x"374" => cos_16 <= x"1B47" ;
        when x"375" => cos_16 <= x"1B16" ;
        when x"376" => cos_16 <= x"1AE5" ;
        when x"377" => cos_16 <= x"1AB4" ;
        when x"378" => cos_16 <= x"1A82" ;
        when x"379" => cos_16 <= x"1A51" ;
        when x"37A" => cos_16 <= x"1A20" ;
        when x"37B" => cos_16 <= x"19EF" ;
        when x"37C" => cos_16 <= x"19BE" ;
        when x"37D" => cos_16 <= x"198C" ;
        when x"37E" => cos_16 <= x"195B" ;
        when x"37F" => cos_16 <= x"192A" ;
        when x"380" => cos_16 <= x"18F9" ;
        when x"381" => cos_16 <= x"18C7" ;
        when x"382" => cos_16 <= x"1896" ;
        when x"383" => cos_16 <= x"1865" ;
        when x"384" => cos_16 <= x"1833" ;
        when x"385" => cos_16 <= x"1802" ;
        when x"386" => cos_16 <= x"17D0" ;
        when x"387" => cos_16 <= x"179F" ;
        when x"388" => cos_16 <= x"176E" ;
        when x"389" => cos_16 <= x"173C" ;
        when x"38A" => cos_16 <= x"170B" ;
        when x"38B" => cos_16 <= x"16D9" ;
        when x"38C" => cos_16 <= x"16A8" ;
        when x"38D" => cos_16 <= x"1676" ;
        when x"38E" => cos_16 <= x"1645" ;
        when x"38F" => cos_16 <= x"1613" ;
        when x"390" => cos_16 <= x"15E2" ;
        when x"391" => cos_16 <= x"15B0" ;
        when x"392" => cos_16 <= x"157F" ;
        when x"393" => cos_16 <= x"154D" ;
        when x"394" => cos_16 <= x"151C" ;
        when x"395" => cos_16 <= x"14EA" ;
        when x"396" => cos_16 <= x"14B9" ;
        when x"397" => cos_16 <= x"1487" ;
        when x"398" => cos_16 <= x"1455" ;
        when x"399" => cos_16 <= x"1424" ;
        when x"39A" => cos_16 <= x"13F2" ;
        when x"39B" => cos_16 <= x"13C0" ;
        when x"39C" => cos_16 <= x"138F" ;
        when x"39D" => cos_16 <= x"135D" ;
        when x"39E" => cos_16 <= x"132B" ;
        when x"39F" => cos_16 <= x"12FA" ;
        when x"3A0" => cos_16 <= x"12C8" ;
        when x"3A1" => cos_16 <= x"1296" ;
        when x"3A2" => cos_16 <= x"1264" ;
        when x"3A3" => cos_16 <= x"1233" ;
        when x"3A4" => cos_16 <= x"1201" ;
        when x"3A5" => cos_16 <= x"11CF" ;
        when x"3A6" => cos_16 <= x"119D" ;
        when x"3A7" => cos_16 <= x"116C" ;
        when x"3A8" => cos_16 <= x"113A" ;
        when x"3A9" => cos_16 <= x"1108" ;
        when x"3AA" => cos_16 <= x"10D6" ;
        when x"3AB" => cos_16 <= x"10A4" ;
        when x"3AC" => cos_16 <= x"1072" ;
        when x"3AD" => cos_16 <= x"1041" ;
        when x"3AE" => cos_16 <= x"100F" ;
        when x"3AF" => cos_16 <= x"0FDD" ;
        when x"3B0" => cos_16 <= x"0FAB" ;
        when x"3B1" => cos_16 <= x"0F79" ;
        when x"3B2" => cos_16 <= x"0F47" ;
        when x"3B3" => cos_16 <= x"0F15" ;
        when x"3B4" => cos_16 <= x"0EE3" ;
        when x"3B5" => cos_16 <= x"0EB1" ;
        when x"3B6" => cos_16 <= x"0E80" ;
        when x"3B7" => cos_16 <= x"0E4E" ;
        when x"3B8" => cos_16 <= x"0E1C" ;
        when x"3B9" => cos_16 <= x"0DEA" ;
        when x"3BA" => cos_16 <= x"0DB8" ;
        when x"3BB" => cos_16 <= x"0D86" ;
        when x"3BC" => cos_16 <= x"0D54" ;
        when x"3BD" => cos_16 <= x"0D22" ;
        when x"3BE" => cos_16 <= x"0CF0" ;
        when x"3BF" => cos_16 <= x"0CBE" ;
        when x"3C0" => cos_16 <= x"0C8C" ;
        when x"3C1" => cos_16 <= x"0C5A" ;
        when x"3C2" => cos_16 <= x"0C28" ;
        when x"3C3" => cos_16 <= x"0BF6" ;
        when x"3C4" => cos_16 <= x"0BC4" ;
        when x"3C5" => cos_16 <= x"0B92" ;
        when x"3C6" => cos_16 <= x"0B5F" ;
        when x"3C7" => cos_16 <= x"0B2D" ;
        when x"3C8" => cos_16 <= x"0AFB" ;
        when x"3C9" => cos_16 <= x"0AC9" ;
        when x"3CA" => cos_16 <= x"0A97" ;
        when x"3CB" => cos_16 <= x"0A65" ;
        when x"3CC" => cos_16 <= x"0A33" ;
        when x"3CD" => cos_16 <= x"0A01" ;
        when x"3CE" => cos_16 <= x"09CF" ;
        when x"3CF" => cos_16 <= x"099D" ;
        when x"3D0" => cos_16 <= x"096A" ;
        when x"3D1" => cos_16 <= x"0938" ;
        when x"3D2" => cos_16 <= x"0906" ;
        when x"3D3" => cos_16 <= x"08D4" ;
        when x"3D4" => cos_16 <= x"08A2" ;
        when x"3D5" => cos_16 <= x"0870" ;
        when x"3D6" => cos_16 <= x"083E" ;
        when x"3D7" => cos_16 <= x"080B" ;
        when x"3D8" => cos_16 <= x"07D9" ;
        when x"3D9" => cos_16 <= x"07A7" ;
        when x"3DA" => cos_16 <= x"0775" ;
        when x"3DB" => cos_16 <= x"0743" ;
        when x"3DC" => cos_16 <= x"0711" ;
        when x"3DD" => cos_16 <= x"06DE" ;
        when x"3DE" => cos_16 <= x"06AC" ;
        when x"3DF" => cos_16 <= x"067A" ;
        when x"3E0" => cos_16 <= x"0648" ;
        when x"3E1" => cos_16 <= x"0616" ;
        when x"3E2" => cos_16 <= x"05E3" ;
        when x"3E3" => cos_16 <= x"05B1" ;
        when x"3E4" => cos_16 <= x"057F" ;
        when x"3E5" => cos_16 <= x"054D" ;
        when x"3E6" => cos_16 <= x"051B" ;
        when x"3E7" => cos_16 <= x"04E8" ;
        when x"3E8" => cos_16 <= x"04B6" ;
        when x"3E9" => cos_16 <= x"0484" ;
        when x"3EA" => cos_16 <= x"0452" ;
        when x"3EB" => cos_16 <= x"041F" ;
        when x"3EC" => cos_16 <= x"03ED" ;
        when x"3ED" => cos_16 <= x"03BB" ;
        when x"3EE" => cos_16 <= x"0389" ;
        when x"3EF" => cos_16 <= x"0356" ;
        when x"3F0" => cos_16 <= x"0324" ;
        when x"3F1" => cos_16 <= x"02F2" ;
        when x"3F2" => cos_16 <= x"02C0" ;
        when x"3F3" => cos_16 <= x"028D" ;
        when x"3F4" => cos_16 <= x"025B" ;
        when x"3F5" => cos_16 <= x"0229" ;
        when x"3F6" => cos_16 <= x"01F7" ;
        when x"3F7" => cos_16 <= x"01C4" ;
        when x"3F8" => cos_16 <= x"0192" ;
        when x"3F9" => cos_16 <= x"0160" ;
        when x"3FA" => cos_16 <= x"012E" ;
        when x"3FB" => cos_16 <= x"00FB" ;
        when x"3FC" => cos_16 <= x"00C9" ;
        when x"3FD" => cos_16 <= x"0097" ;
        when x"3FE" => cos_16 <= x"0065" ;
        when x"3FF" => cos_16 <= x"0032" ;
        when x"400" => cos_16 <= x"0000" ;
        when x"401" => cos_16 <= x"FFCE" ;
        when x"402" => cos_16 <= x"FF9B" ;
        when x"403" => cos_16 <= x"FF69" ;
        when x"404" => cos_16 <= x"FF37" ;
        when x"405" => cos_16 <= x"FF05" ;
        when x"406" => cos_16 <= x"FED2" ;
        when x"407" => cos_16 <= x"FEA0" ;
        when x"408" => cos_16 <= x"FE6E" ;
        when x"409" => cos_16 <= x"FE3C" ;
        when x"40A" => cos_16 <= x"FE09" ;
        when x"40B" => cos_16 <= x"FDD7" ;
        when x"40C" => cos_16 <= x"FDA5" ;
        when x"40D" => cos_16 <= x"FD73" ;
        when x"40E" => cos_16 <= x"FD40" ;
        when x"40F" => cos_16 <= x"FD0E" ;
        when x"410" => cos_16 <= x"FCDC" ;
        when x"411" => cos_16 <= x"FCAA" ;
        when x"412" => cos_16 <= x"FC77" ;
        when x"413" => cos_16 <= x"FC45" ;
        when x"414" => cos_16 <= x"FC13" ;
        when x"415" => cos_16 <= x"FBE1" ;
        when x"416" => cos_16 <= x"FBAE" ;
        when x"417" => cos_16 <= x"FB7C" ;
        when x"418" => cos_16 <= x"FB4A" ;
        when x"419" => cos_16 <= x"FB18" ;
        when x"41A" => cos_16 <= x"FAE5" ;
        when x"41B" => cos_16 <= x"FAB3" ;
        when x"41C" => cos_16 <= x"FA81" ;
        when x"41D" => cos_16 <= x"FA4F" ;
        when x"41E" => cos_16 <= x"FA1D" ;
        when x"41F" => cos_16 <= x"F9EA" ;
        when x"420" => cos_16 <= x"F9B8" ;
        when x"421" => cos_16 <= x"F986" ;
        when x"422" => cos_16 <= x"F954" ;
        when x"423" => cos_16 <= x"F922" ;
        when x"424" => cos_16 <= x"F8EF" ;
        when x"425" => cos_16 <= x"F8BD" ;
        when x"426" => cos_16 <= x"F88B" ;
        when x"427" => cos_16 <= x"F859" ;
        when x"428" => cos_16 <= x"F827" ;
        when x"429" => cos_16 <= x"F7F5" ;
        when x"42A" => cos_16 <= x"F7C2" ;
        when x"42B" => cos_16 <= x"F790" ;
        when x"42C" => cos_16 <= x"F75E" ;
        when x"42D" => cos_16 <= x"F72C" ;
        when x"42E" => cos_16 <= x"F6FA" ;
        when x"42F" => cos_16 <= x"F6C8" ;
        when x"430" => cos_16 <= x"F696" ;
        when x"431" => cos_16 <= x"F663" ;
        when x"432" => cos_16 <= x"F631" ;
        when x"433" => cos_16 <= x"F5FF" ;
        when x"434" => cos_16 <= x"F5CD" ;
        when x"435" => cos_16 <= x"F59B" ;
        when x"436" => cos_16 <= x"F569" ;
        when x"437" => cos_16 <= x"F537" ;
        when x"438" => cos_16 <= x"F505" ;
        when x"439" => cos_16 <= x"F4D3" ;
        when x"43A" => cos_16 <= x"F4A1" ;
        when x"43B" => cos_16 <= x"F46E" ;
        when x"43C" => cos_16 <= x"F43C" ;
        when x"43D" => cos_16 <= x"F40A" ;
        when x"43E" => cos_16 <= x"F3D8" ;
        when x"43F" => cos_16 <= x"F3A6" ;
        when x"440" => cos_16 <= x"F374" ;
        when x"441" => cos_16 <= x"F342" ;
        when x"442" => cos_16 <= x"F310" ;
        when x"443" => cos_16 <= x"F2DE" ;
        when x"444" => cos_16 <= x"F2AC" ;
        when x"445" => cos_16 <= x"F27A" ;
        when x"446" => cos_16 <= x"F248" ;
        when x"447" => cos_16 <= x"F216" ;
        when x"448" => cos_16 <= x"F1E4" ;
        when x"449" => cos_16 <= x"F1B2" ;
        when x"44A" => cos_16 <= x"F180" ;
        when x"44B" => cos_16 <= x"F14F" ;
        when x"44C" => cos_16 <= x"F11D" ;
        when x"44D" => cos_16 <= x"F0EB" ;
        when x"44E" => cos_16 <= x"F0B9" ;
        when x"44F" => cos_16 <= x"F087" ;
        when x"450" => cos_16 <= x"F055" ;
        when x"451" => cos_16 <= x"F023" ;
        when x"452" => cos_16 <= x"EFF1" ;
        when x"453" => cos_16 <= x"EFBF" ;
        when x"454" => cos_16 <= x"EF8E" ;
        when x"455" => cos_16 <= x"EF5C" ;
        when x"456" => cos_16 <= x"EF2A" ;
        when x"457" => cos_16 <= x"EEF8" ;
        when x"458" => cos_16 <= x"EEC6" ;
        when x"459" => cos_16 <= x"EE94" ;
        when x"45A" => cos_16 <= x"EE63" ;
        when x"45B" => cos_16 <= x"EE31" ;
        when x"45C" => cos_16 <= x"EDFF" ;
        when x"45D" => cos_16 <= x"EDCD" ;
        when x"45E" => cos_16 <= x"ED9C" ;
        when x"45F" => cos_16 <= x"ED6A" ;
        when x"460" => cos_16 <= x"ED38" ;
        when x"461" => cos_16 <= x"ED06" ;
        when x"462" => cos_16 <= x"ECD5" ;
        when x"463" => cos_16 <= x"ECA3" ;
        when x"464" => cos_16 <= x"EC71" ;
        when x"465" => cos_16 <= x"EC40" ;
        when x"466" => cos_16 <= x"EC0E" ;
        when x"467" => cos_16 <= x"EBDC" ;
        when x"468" => cos_16 <= x"EBAB" ;
        when x"469" => cos_16 <= x"EB79" ;
        when x"46A" => cos_16 <= x"EB47" ;
        when x"46B" => cos_16 <= x"EB16" ;
        when x"46C" => cos_16 <= x"EAE4" ;
        when x"46D" => cos_16 <= x"EAB3" ;
        when x"46E" => cos_16 <= x"EA81" ;
        when x"46F" => cos_16 <= x"EA50" ;
        when x"470" => cos_16 <= x"EA1E" ;
        when x"471" => cos_16 <= x"E9ED" ;
        when x"472" => cos_16 <= x"E9BB" ;
        when x"473" => cos_16 <= x"E98A" ;
        when x"474" => cos_16 <= x"E958" ;
        when x"475" => cos_16 <= x"E927" ;
        when x"476" => cos_16 <= x"E8F5" ;
        when x"477" => cos_16 <= x"E8C4" ;
        when x"478" => cos_16 <= x"E892" ;
        when x"479" => cos_16 <= x"E861" ;
        when x"47A" => cos_16 <= x"E830" ;
        when x"47B" => cos_16 <= x"E7FE" ;
        when x"47C" => cos_16 <= x"E7CD" ;
        when x"47D" => cos_16 <= x"E79B" ;
        when x"47E" => cos_16 <= x"E76A" ;
        when x"47F" => cos_16 <= x"E739" ;
        when x"480" => cos_16 <= x"E707" ;
        when x"481" => cos_16 <= x"E6D6" ;
        when x"482" => cos_16 <= x"E6A5" ;
        when x"483" => cos_16 <= x"E674" ;
        when x"484" => cos_16 <= x"E642" ;
        when x"485" => cos_16 <= x"E611" ;
        when x"486" => cos_16 <= x"E5E0" ;
        when x"487" => cos_16 <= x"E5AF" ;
        when x"488" => cos_16 <= x"E57E" ;
        when x"489" => cos_16 <= x"E54C" ;
        when x"48A" => cos_16 <= x"E51B" ;
        when x"48B" => cos_16 <= x"E4EA" ;
        when x"48C" => cos_16 <= x"E4B9" ;
        when x"48D" => cos_16 <= x"E488" ;
        when x"48E" => cos_16 <= x"E457" ;
        when x"48F" => cos_16 <= x"E426" ;
        when x"490" => cos_16 <= x"E3F5" ;
        when x"491" => cos_16 <= x"E3C4" ;
        when x"492" => cos_16 <= x"E393" ;
        when x"493" => cos_16 <= x"E362" ;
        when x"494" => cos_16 <= x"E331" ;
        when x"495" => cos_16 <= x"E300" ;
        when x"496" => cos_16 <= x"E2CF" ;
        when x"497" => cos_16 <= x"E29E" ;
        when x"498" => cos_16 <= x"E26D" ;
        when x"499" => cos_16 <= x"E23C" ;
        when x"49A" => cos_16 <= x"E20B" ;
        when x"49B" => cos_16 <= x"E1DA" ;
        when x"49C" => cos_16 <= x"E1A9" ;
        when x"49D" => cos_16 <= x"E179" ;
        when x"49E" => cos_16 <= x"E148" ;
        when x"49F" => cos_16 <= x"E117" ;
        when x"4A0" => cos_16 <= x"E0E6" ;
        when x"4A1" => cos_16 <= x"E0B6" ;
        when x"4A2" => cos_16 <= x"E085" ;
        when x"4A3" => cos_16 <= x"E054" ;
        when x"4A4" => cos_16 <= x"E023" ;
        when x"4A5" => cos_16 <= x"DFF3" ;
        when x"4A6" => cos_16 <= x"DFC2" ;
        when x"4A7" => cos_16 <= x"DF91" ;
        when x"4A8" => cos_16 <= x"DF61" ;
        when x"4A9" => cos_16 <= x"DF30" ;
        when x"4AA" => cos_16 <= x"DF00" ;
        when x"4AB" => cos_16 <= x"DECF" ;
        when x"4AC" => cos_16 <= x"DE9F" ;
        when x"4AD" => cos_16 <= x"DE6E" ;
        when x"4AE" => cos_16 <= x"DE3E" ;
        when x"4AF" => cos_16 <= x"DE0D" ;
        when x"4B0" => cos_16 <= x"DDDD" ;
        when x"4B1" => cos_16 <= x"DDAC" ;
        when x"4B2" => cos_16 <= x"DD7C" ;
        when x"4B3" => cos_16 <= x"DD4B" ;
        when x"4B4" => cos_16 <= x"DD1B" ;
        when x"4B5" => cos_16 <= x"DCEB" ;
        when x"4B6" => cos_16 <= x"DCBA" ;
        when x"4B7" => cos_16 <= x"DC8A" ;
        when x"4B8" => cos_16 <= x"DC5A" ;
        when x"4B9" => cos_16 <= x"DC29" ;
        when x"4BA" => cos_16 <= x"DBF9" ;
        when x"4BB" => cos_16 <= x"DBC9" ;
        when x"4BC" => cos_16 <= x"DB99" ;
        when x"4BD" => cos_16 <= x"DB69" ;
        when x"4BE" => cos_16 <= x"DB38" ;
        when x"4BF" => cos_16 <= x"DB08" ;
        when x"4C0" => cos_16 <= x"DAD8" ;
        when x"4C1" => cos_16 <= x"DAA8" ;
        when x"4C2" => cos_16 <= x"DA78" ;
        when x"4C3" => cos_16 <= x"DA48" ;
        when x"4C4" => cos_16 <= x"DA18" ;
        when x"4C5" => cos_16 <= x"D9E8" ;
        when x"4C6" => cos_16 <= x"D9B8" ;
        when x"4C7" => cos_16 <= x"D988" ;
        when x"4C8" => cos_16 <= x"D958" ;
        when x"4C9" => cos_16 <= x"D928" ;
        when x"4CA" => cos_16 <= x"D8F8" ;
        when x"4CB" => cos_16 <= x"D8C9" ;
        when x"4CC" => cos_16 <= x"D899" ;
        when x"4CD" => cos_16 <= x"D869" ;
        when x"4CE" => cos_16 <= x"D839" ;
        when x"4CF" => cos_16 <= x"D809" ;
        when x"4D0" => cos_16 <= x"D7DA" ;
        when x"4D1" => cos_16 <= x"D7AA" ;
        when x"4D2" => cos_16 <= x"D77A" ;
        when x"4D3" => cos_16 <= x"D74B" ;
        when x"4D4" => cos_16 <= x"D71B" ;
        when x"4D5" => cos_16 <= x"D6EB" ;
        when x"4D6" => cos_16 <= x"D6BC" ;
        when x"4D7" => cos_16 <= x"D68C" ;
        when x"4D8" => cos_16 <= x"D65D" ;
        when x"4D9" => cos_16 <= x"D62D" ;
        when x"4DA" => cos_16 <= x"D5FE" ;
        when x"4DB" => cos_16 <= x"D5CE" ;
        when x"4DC" => cos_16 <= x"D59F" ;
        when x"4DD" => cos_16 <= x"D56F" ;
        when x"4DE" => cos_16 <= x"D540" ;
        when x"4DF" => cos_16 <= x"D510" ;
        when x"4E0" => cos_16 <= x"D4E1" ;
        when x"4E1" => cos_16 <= x"D4B2" ;
        when x"4E2" => cos_16 <= x"D483" ;
        when x"4E3" => cos_16 <= x"D453" ;
        when x"4E4" => cos_16 <= x"D424" ;
        when x"4E5" => cos_16 <= x"D3F5" ;
        when x"4E6" => cos_16 <= x"D3C6" ;
        when x"4E7" => cos_16 <= x"D396" ;
        when x"4E8" => cos_16 <= x"D367" ;
        when x"4E9" => cos_16 <= x"D338" ;
        when x"4EA" => cos_16 <= x"D309" ;
        when x"4EB" => cos_16 <= x"D2DA" ;
        when x"4EC" => cos_16 <= x"D2AB" ;
        when x"4ED" => cos_16 <= x"D27C" ;
        when x"4EE" => cos_16 <= x"D24D" ;
        when x"4EF" => cos_16 <= x"D21E" ;
        when x"4F0" => cos_16 <= x"D1EF" ;
        when x"4F1" => cos_16 <= x"D1C0" ;
        when x"4F2" => cos_16 <= x"D192" ;
        when x"4F3" => cos_16 <= x"D163" ;
        when x"4F4" => cos_16 <= x"D134" ;
        when x"4F5" => cos_16 <= x"D105" ;
        when x"4F6" => cos_16 <= x"D0D6" ;
        when x"4F7" => cos_16 <= x"D0A8" ;
        when x"4F8" => cos_16 <= x"D079" ;
        when x"4F9" => cos_16 <= x"D04A" ;
        when x"4FA" => cos_16 <= x"D01C" ;
        when x"4FB" => cos_16 <= x"CFED" ;
        when x"4FC" => cos_16 <= x"CFBF" ;
        when x"4FD" => cos_16 <= x"CF90" ;
        when x"4FE" => cos_16 <= x"CF62" ;
        when x"4FF" => cos_16 <= x"CF33" ;
        when x"500" => cos_16 <= x"CF05" ;
        when x"501" => cos_16 <= x"CED6" ;
        when x"502" => cos_16 <= x"CEA8" ;
        when x"503" => cos_16 <= x"CE79" ;
        when x"504" => cos_16 <= x"CE4B" ;
        when x"505" => cos_16 <= x"CE1D" ;
        when x"506" => cos_16 <= x"CDEF" ;
        when x"507" => cos_16 <= x"CDC0" ;
        when x"508" => cos_16 <= x"CD92" ;
        when x"509" => cos_16 <= x"CD64" ;
        when x"50A" => cos_16 <= x"CD36" ;
        when x"50B" => cos_16 <= x"CD08" ;
        when x"50C" => cos_16 <= x"CCDA" ;
        when x"50D" => cos_16 <= x"CCAB" ;
        when x"50E" => cos_16 <= x"CC7D" ;
        when x"50F" => cos_16 <= x"CC4F" ;
        when x"510" => cos_16 <= x"CC21" ;
        when x"511" => cos_16 <= x"CBF4" ;
        when x"512" => cos_16 <= x"CBC6" ;
        when x"513" => cos_16 <= x"CB98" ;
        when x"514" => cos_16 <= x"CB6A" ;
        when x"515" => cos_16 <= x"CB3C" ;
        when x"516" => cos_16 <= x"CB0E" ;
        when x"517" => cos_16 <= x"CAE1" ;
        when x"518" => cos_16 <= x"CAB3" ;
        when x"519" => cos_16 <= x"CA85" ;
        when x"51A" => cos_16 <= x"CA58" ;
        when x"51B" => cos_16 <= x"CA2A" ;
        when x"51C" => cos_16 <= x"C9FC" ;
        when x"51D" => cos_16 <= x"C9CF" ;
        when x"51E" => cos_16 <= x"C9A1" ;
        when x"51F" => cos_16 <= x"C974" ;
        when x"520" => cos_16 <= x"C946" ;
        when x"521" => cos_16 <= x"C919" ;
        when x"522" => cos_16 <= x"C8EB" ;
        when x"523" => cos_16 <= x"C8BE" ;
        when x"524" => cos_16 <= x"C891" ;
        when x"525" => cos_16 <= x"C864" ;
        when x"526" => cos_16 <= x"C836" ;
        when x"527" => cos_16 <= x"C809" ;
        when x"528" => cos_16 <= x"C7DC" ;
        when x"529" => cos_16 <= x"C7AF" ;
        when x"52A" => cos_16 <= x"C782" ;
        when x"52B" => cos_16 <= x"C755" ;
        when x"52C" => cos_16 <= x"C727" ;
        when x"52D" => cos_16 <= x"C6FA" ;
        when x"52E" => cos_16 <= x"C6CD" ;
        when x"52F" => cos_16 <= x"C6A0" ;
        when x"530" => cos_16 <= x"C674" ;
        when x"531" => cos_16 <= x"C647" ;
        when x"532" => cos_16 <= x"C61A" ;
        when x"533" => cos_16 <= x"C5ED" ;
        when x"534" => cos_16 <= x"C5C0" ;
        when x"535" => cos_16 <= x"C594" ;
        when x"536" => cos_16 <= x"C567" ;
        when x"537" => cos_16 <= x"C53A" ;
        when x"538" => cos_16 <= x"C50E" ;
        when x"539" => cos_16 <= x"C4E1" ;
        when x"53A" => cos_16 <= x"C4B4" ;
        when x"53B" => cos_16 <= x"C488" ;
        when x"53C" => cos_16 <= x"C45B" ;
        when x"53D" => cos_16 <= x"C42F" ;
        when x"53E" => cos_16 <= x"C402" ;
        when x"53F" => cos_16 <= x"C3D6" ;
        when x"540" => cos_16 <= x"C3AA" ;
        when x"541" => cos_16 <= x"C37D" ;
        when x"542" => cos_16 <= x"C351" ;
        when x"543" => cos_16 <= x"C325" ;
        when x"544" => cos_16 <= x"C2F9" ;
        when x"545" => cos_16 <= x"C2CD" ;
        when x"546" => cos_16 <= x"C2A0" ;
        when x"547" => cos_16 <= x"C274" ;
        when x"548" => cos_16 <= x"C248" ;
        when x"549" => cos_16 <= x"C21C" ;
        when x"54A" => cos_16 <= x"C1F0" ;
        when x"54B" => cos_16 <= x"C1C4" ;
        when x"54C" => cos_16 <= x"C198" ;
        when x"54D" => cos_16 <= x"C16D" ;
        when x"54E" => cos_16 <= x"C141" ;
        when x"54F" => cos_16 <= x"C115" ;
        when x"550" => cos_16 <= x"C0E9" ;
        when x"551" => cos_16 <= x"C0BD" ;
        when x"552" => cos_16 <= x"C092" ;
        when x"553" => cos_16 <= x"C066" ;
        when x"554" => cos_16 <= x"C03B" ;
        when x"555" => cos_16 <= x"C00F" ;
        when x"556" => cos_16 <= x"BFE3" ;
        when x"557" => cos_16 <= x"BFB8" ;
        when x"558" => cos_16 <= x"BF8D" ;
        when x"559" => cos_16 <= x"BF61" ;
        when x"55A" => cos_16 <= x"BF36" ;
        when x"55B" => cos_16 <= x"BF0A" ;
        when x"55C" => cos_16 <= x"BEDF" ;
        when x"55D" => cos_16 <= x"BEB4" ;
        when x"55E" => cos_16 <= x"BE89" ;
        when x"55F" => cos_16 <= x"BE5E" ;
        when x"560" => cos_16 <= x"BE32" ;
        when x"561" => cos_16 <= x"BE07" ;
        when x"562" => cos_16 <= x"BDDC" ;
        when x"563" => cos_16 <= x"BDB1" ;
        when x"564" => cos_16 <= x"BD86" ;
        when x"565" => cos_16 <= x"BD5B" ;
        when x"566" => cos_16 <= x"BD30" ;
        when x"567" => cos_16 <= x"BD06" ;
        when x"568" => cos_16 <= x"BCDB" ;
        when x"569" => cos_16 <= x"BCB0" ;
        when x"56A" => cos_16 <= x"BC85" ;
        when x"56B" => cos_16 <= x"BC5B" ;
        when x"56C" => cos_16 <= x"BC30" ;
        when x"56D" => cos_16 <= x"BC05" ;
        when x"56E" => cos_16 <= x"BBDB" ;
        when x"56F" => cos_16 <= x"BBB0" ;
        when x"570" => cos_16 <= x"BB86" ;
        when x"571" => cos_16 <= x"BB5B" ;
        when x"572" => cos_16 <= x"BB31" ;
        when x"573" => cos_16 <= x"BB07" ;
        when x"574" => cos_16 <= x"BADC" ;
        when x"575" => cos_16 <= x"BAB2" ;
        when x"576" => cos_16 <= x"BA88" ;
        when x"577" => cos_16 <= x"BA5D" ;
        when x"578" => cos_16 <= x"BA33" ;
        when x"579" => cos_16 <= x"BA09" ;
        when x"57A" => cos_16 <= x"B9DF" ;
        when x"57B" => cos_16 <= x"B9B5" ;
        when x"57C" => cos_16 <= x"B98B" ;
        when x"57D" => cos_16 <= x"B961" ;
        when x"57E" => cos_16 <= x"B937" ;
        when x"57F" => cos_16 <= x"B90D" ;
        when x"580" => cos_16 <= x"B8E4" ;
        when x"581" => cos_16 <= x"B8BA" ;
        when x"582" => cos_16 <= x"B890" ;
        when x"583" => cos_16 <= x"B866" ;
        when x"584" => cos_16 <= x"B83D" ;
        when x"585" => cos_16 <= x"B813" ;
        when x"586" => cos_16 <= x"B7EA" ;
        when x"587" => cos_16 <= x"B7C0" ;
        when x"588" => cos_16 <= x"B797" ;
        when x"589" => cos_16 <= x"B76D" ;
        when x"58A" => cos_16 <= x"B744" ;
        when x"58B" => cos_16 <= x"B71B" ;
        when x"58C" => cos_16 <= x"B6F1" ;
        when x"58D" => cos_16 <= x"B6C8" ;
        when x"58E" => cos_16 <= x"B69F" ;
        when x"58F" => cos_16 <= x"B676" ;
        when x"590" => cos_16 <= x"B64C" ;
        when x"591" => cos_16 <= x"B623" ;
        when x"592" => cos_16 <= x"B5FA" ;
        when x"593" => cos_16 <= x"B5D1" ;
        when x"594" => cos_16 <= x"B5A8" ;
        when x"595" => cos_16 <= x"B580" ;
        when x"596" => cos_16 <= x"B557" ;
        when x"597" => cos_16 <= x"B52E" ;
        when x"598" => cos_16 <= x"B505" ;
        when x"599" => cos_16 <= x"B4DC" ;
        when x"59A" => cos_16 <= x"B4B4" ;
        when x"59B" => cos_16 <= x"B48B" ;
        when x"59C" => cos_16 <= x"B463" ;
        when x"59D" => cos_16 <= x"B43A" ;
        when x"59E" => cos_16 <= x"B412" ;
        when x"59F" => cos_16 <= x"B3E9" ;
        when x"5A0" => cos_16 <= x"B3C1" ;
        when x"5A1" => cos_16 <= x"B398" ;
        when x"5A2" => cos_16 <= x"B370" ;
        when x"5A3" => cos_16 <= x"B348" ;
        when x"5A4" => cos_16 <= x"B320" ;
        when x"5A5" => cos_16 <= x"B2F7" ;
        when x"5A6" => cos_16 <= x"B2CF" ;
        when x"5A7" => cos_16 <= x"B2A7" ;
        when x"5A8" => cos_16 <= x"B27F" ;
        when x"5A9" => cos_16 <= x"B257" ;
        when x"5AA" => cos_16 <= x"B22F" ;
        when x"5AB" => cos_16 <= x"B207" ;
        when x"5AC" => cos_16 <= x"B1E0" ;
        when x"5AD" => cos_16 <= x"B1B8" ;
        when x"5AE" => cos_16 <= x"B190" ;
        when x"5AF" => cos_16 <= x"B168" ;
        when x"5B0" => cos_16 <= x"B141" ;
        when x"5B1" => cos_16 <= x"B119" ;
        when x"5B2" => cos_16 <= x"B0F2" ;
        when x"5B3" => cos_16 <= x"B0CA" ;
        when x"5B4" => cos_16 <= x"B0A3" ;
        when x"5B5" => cos_16 <= x"B07B" ;
        when x"5B6" => cos_16 <= x"B054" ;
        when x"5B7" => cos_16 <= x"B02C" ;
        when x"5B8" => cos_16 <= x"B005" ;
        when x"5B9" => cos_16 <= x"AFDE" ;
        when x"5BA" => cos_16 <= x"AFB7" ;
        when x"5BB" => cos_16 <= x"AF90" ;
        when x"5BC" => cos_16 <= x"AF69" ;
        when x"5BD" => cos_16 <= x"AF42" ;
        when x"5BE" => cos_16 <= x"AF1B" ;
        when x"5BF" => cos_16 <= x"AEF4" ;
        when x"5C0" => cos_16 <= x"AECD" ;
        when x"5C1" => cos_16 <= x"AEA6" ;
        when x"5C2" => cos_16 <= x"AE7F" ;
        when x"5C3" => cos_16 <= x"AE58" ;
        when x"5C4" => cos_16 <= x"AE32" ;
        when x"5C5" => cos_16 <= x"AE0B" ;
        when x"5C6" => cos_16 <= x"ADE5" ;
        when x"5C7" => cos_16 <= x"ADBE" ;
        when x"5C8" => cos_16 <= x"AD98" ;
        when x"5C9" => cos_16 <= x"AD71" ;
        when x"5CA" => cos_16 <= x"AD4B" ;
        when x"5CB" => cos_16 <= x"AD24" ;
        when x"5CC" => cos_16 <= x"ACFE" ;
        when x"5CD" => cos_16 <= x"ACD8" ;
        when x"5CE" => cos_16 <= x"ACB2" ;
        when x"5CF" => cos_16 <= x"AC8C" ;
        when x"5D0" => cos_16 <= x"AC65" ;
        when x"5D1" => cos_16 <= x"AC3F" ;
        when x"5D2" => cos_16 <= x"AC19" ;
        when x"5D3" => cos_16 <= x"ABF4" ;
        when x"5D4" => cos_16 <= x"ABCE" ;
        when x"5D5" => cos_16 <= x"ABA8" ;
        when x"5D6" => cos_16 <= x"AB82" ;
        when x"5D7" => cos_16 <= x"AB5C" ;
        when x"5D8" => cos_16 <= x"AB37" ;
        when x"5D9" => cos_16 <= x"AB11" ;
        when x"5DA" => cos_16 <= x"AAEB" ;
        when x"5DB" => cos_16 <= x"AAC6" ;
        when x"5DC" => cos_16 <= x"AAA0" ;
        when x"5DD" => cos_16 <= x"AA7B" ;
        when x"5DE" => cos_16 <= x"AA56" ;
        when x"5DF" => cos_16 <= x"AA30" ;
        when x"5E0" => cos_16 <= x"AA0B" ;
        when x"5E1" => cos_16 <= x"A9E6" ;
        when x"5E2" => cos_16 <= x"A9C1" ;
        when x"5E3" => cos_16 <= x"A99C" ;
        when x"5E4" => cos_16 <= x"A976" ;
        when x"5E5" => cos_16 <= x"A951" ;
        when x"5E6" => cos_16 <= x"A92D" ;
        when x"5E7" => cos_16 <= x"A908" ;
        when x"5E8" => cos_16 <= x"A8E3" ;
        when x"5E9" => cos_16 <= x"A8BE" ;
        when x"5EA" => cos_16 <= x"A899" ;
        when x"5EB" => cos_16 <= x"A875" ;
        when x"5EC" => cos_16 <= x"A850" ;
        when x"5ED" => cos_16 <= x"A82B" ;
        when x"5EE" => cos_16 <= x"A807" ;
        when x"5EF" => cos_16 <= x"A7E2" ;
        when x"5F0" => cos_16 <= x"A7BE" ;
        when x"5F1" => cos_16 <= x"A799" ;
        when x"5F2" => cos_16 <= x"A775" ;
        when x"5F3" => cos_16 <= x"A751" ;
        when x"5F4" => cos_16 <= x"A72D" ;
        when x"5F5" => cos_16 <= x"A708" ;
        when x"5F6" => cos_16 <= x"A6E4" ;
        when x"5F7" => cos_16 <= x"A6C0" ;
        when x"5F8" => cos_16 <= x"A69C" ;
        when x"5F9" => cos_16 <= x"A678" ;
        when x"5FA" => cos_16 <= x"A654" ;
        when x"5FB" => cos_16 <= x"A631" ;
        when x"5FC" => cos_16 <= x"A60D" ;
        when x"5FD" => cos_16 <= x"A5E9" ;
        when x"5FE" => cos_16 <= x"A5C5" ;
        when x"5FF" => cos_16 <= x"A5A2" ;
        when x"600" => cos_16 <= x"A57E" ;
        when x"601" => cos_16 <= x"A55B" ;
        when x"602" => cos_16 <= x"A537" ;
        when x"603" => cos_16 <= x"A514" ;
        when x"604" => cos_16 <= x"A4F1" ;
        when x"605" => cos_16 <= x"A4CD" ;
        when x"606" => cos_16 <= x"A4AA" ;
        when x"607" => cos_16 <= x"A487" ;
        when x"608" => cos_16 <= x"A464" ;
        when x"609" => cos_16 <= x"A441" ;
        when x"60A" => cos_16 <= x"A41E" ;
        when x"60B" => cos_16 <= x"A3FB" ;
        when x"60C" => cos_16 <= x"A3D8" ;
        when x"60D" => cos_16 <= x"A3B5" ;
        when x"60E" => cos_16 <= x"A392" ;
        when x"60F" => cos_16 <= x"A36F" ;
        when x"610" => cos_16 <= x"A34D" ;
        when x"611" => cos_16 <= x"A32A" ;
        when x"612" => cos_16 <= x"A307" ;
        when x"613" => cos_16 <= x"A2E5" ;
        when x"614" => cos_16 <= x"A2C2" ;
        when x"615" => cos_16 <= x"A2A0" ;
        when x"616" => cos_16 <= x"A27E" ;
        when x"617" => cos_16 <= x"A25B" ;
        when x"618" => cos_16 <= x"A239" ;
        when x"619" => cos_16 <= x"A217" ;
        when x"61A" => cos_16 <= x"A1F5" ;
        when x"61B" => cos_16 <= x"A1D3" ;
        when x"61C" => cos_16 <= x"A1B1" ;
        when x"61D" => cos_16 <= x"A18F" ;
        when x"61E" => cos_16 <= x"A16D" ;
        when x"61F" => cos_16 <= x"A14B" ;
        when x"620" => cos_16 <= x"A129" ;
        when x"621" => cos_16 <= x"A108" ;
        when x"622" => cos_16 <= x"A0E6" ;
        when x"623" => cos_16 <= x"A0C4" ;
        when x"624" => cos_16 <= x"A0A3" ;
        when x"625" => cos_16 <= x"A081" ;
        when x"626" => cos_16 <= x"A060" ;
        when x"627" => cos_16 <= x"A03E" ;
        when x"628" => cos_16 <= x"A01D" ;
        when x"629" => cos_16 <= x"9FFC" ;
        when x"62A" => cos_16 <= x"9FDB" ;
        when x"62B" => cos_16 <= x"9FB9" ;
        when x"62C" => cos_16 <= x"9F98" ;
        when x"62D" => cos_16 <= x"9F77" ;
        when x"62E" => cos_16 <= x"9F56" ;
        when x"62F" => cos_16 <= x"9F35" ;
        when x"630" => cos_16 <= x"9F15" ;
        when x"631" => cos_16 <= x"9EF4" ;
        when x"632" => cos_16 <= x"9ED3" ;
        when x"633" => cos_16 <= x"9EB2" ;
        when x"634" => cos_16 <= x"9E92" ;
        when x"635" => cos_16 <= x"9E71" ;
        when x"636" => cos_16 <= x"9E51" ;
        when x"637" => cos_16 <= x"9E30" ;
        when x"638" => cos_16 <= x"9E10" ;
        when x"639" => cos_16 <= x"9DEF" ;
        when x"63A" => cos_16 <= x"9DCF" ;
        when x"63B" => cos_16 <= x"9DAF" ;
        when x"63C" => cos_16 <= x"9D8F" ;
        when x"63D" => cos_16 <= x"9D6F" ;
        when x"63E" => cos_16 <= x"9D4F" ;
        when x"63F" => cos_16 <= x"9D2F" ;
        when x"640" => cos_16 <= x"9D0F" ;
        when x"641" => cos_16 <= x"9CEF" ;
        when x"642" => cos_16 <= x"9CCF" ;
        when x"643" => cos_16 <= x"9CAF" ;
        when x"644" => cos_16 <= x"9C90" ;
        when x"645" => cos_16 <= x"9C70" ;
        when x"646" => cos_16 <= x"9C51" ;
        when x"647" => cos_16 <= x"9C31" ;
        when x"648" => cos_16 <= x"9C12" ;
        when x"649" => cos_16 <= x"9BF2" ;
        when x"64A" => cos_16 <= x"9BD3" ;
        when x"64B" => cos_16 <= x"9BB4" ;
        when x"64C" => cos_16 <= x"9B94" ;
        when x"64D" => cos_16 <= x"9B75" ;
        when x"64E" => cos_16 <= x"9B56" ;
        when x"64F" => cos_16 <= x"9B37" ;
        when x"650" => cos_16 <= x"9B18" ;
        when x"651" => cos_16 <= x"9AF9" ;
        when x"652" => cos_16 <= x"9ADB" ;
        when x"653" => cos_16 <= x"9ABC" ;
        when x"654" => cos_16 <= x"9A9D" ;
        when x"655" => cos_16 <= x"9A7E" ;
        when x"656" => cos_16 <= x"9A60" ;
        when x"657" => cos_16 <= x"9A41" ;
        when x"658" => cos_16 <= x"9A23" ;
        when x"659" => cos_16 <= x"9A04" ;
        when x"65A" => cos_16 <= x"99E6" ;
        when x"65B" => cos_16 <= x"99C8" ;
        when x"65C" => cos_16 <= x"99AA" ;
        when x"65D" => cos_16 <= x"998B" ;
        when x"65E" => cos_16 <= x"996D" ;
        when x"65F" => cos_16 <= x"994F" ;
        when x"660" => cos_16 <= x"9931" ;
        when x"661" => cos_16 <= x"9913" ;
        when x"662" => cos_16 <= x"98F6" ;
        when x"663" => cos_16 <= x"98D8" ;
        when x"664" => cos_16 <= x"98BA" ;
        when x"665" => cos_16 <= x"989C" ;
        when x"666" => cos_16 <= x"987F" ;
        when x"667" => cos_16 <= x"9861" ;
        when x"668" => cos_16 <= x"9844" ;
        when x"669" => cos_16 <= x"9826" ;
        when x"66A" => cos_16 <= x"9809" ;
        when x"66B" => cos_16 <= x"97EC" ;
        when x"66C" => cos_16 <= x"97CE" ;
        when x"66D" => cos_16 <= x"97B1" ;
        when x"66E" => cos_16 <= x"9794" ;
        when x"66F" => cos_16 <= x"9777" ;
        when x"670" => cos_16 <= x"975A" ;
        when x"671" => cos_16 <= x"973D" ;
        when x"672" => cos_16 <= x"9720" ;
        when x"673" => cos_16 <= x"9704" ;
        when x"674" => cos_16 <= x"96E7" ;
        when x"675" => cos_16 <= x"96CA" ;
        when x"676" => cos_16 <= x"96AE" ;
        when x"677" => cos_16 <= x"9691" ;
        when x"678" => cos_16 <= x"9675" ;
        when x"679" => cos_16 <= x"9658" ;
        when x"67A" => cos_16 <= x"963C" ;
        when x"67B" => cos_16 <= x"9620" ;
        when x"67C" => cos_16 <= x"9603" ;
        when x"67D" => cos_16 <= x"95E7" ;
        when x"67E" => cos_16 <= x"95CB" ;
        when x"67F" => cos_16 <= x"95AF" ;
        when x"680" => cos_16 <= x"9593" ;
        when x"681" => cos_16 <= x"9577" ;
        when x"682" => cos_16 <= x"955C" ;
        when x"683" => cos_16 <= x"9540" ;
        when x"684" => cos_16 <= x"9524" ;
        when x"685" => cos_16 <= x"9508" ;
        when x"686" => cos_16 <= x"94ED" ;
        when x"687" => cos_16 <= x"94D1" ;
        when x"688" => cos_16 <= x"94B6" ;
        when x"689" => cos_16 <= x"949B" ;
        when x"68A" => cos_16 <= x"947F" ;
        when x"68B" => cos_16 <= x"9464" ;
        when x"68C" => cos_16 <= x"9449" ;
        when x"68D" => cos_16 <= x"942E" ;
        when x"68E" => cos_16 <= x"9413" ;
        when x"68F" => cos_16 <= x"93F8" ;
        when x"690" => cos_16 <= x"93DD" ;
        when x"691" => cos_16 <= x"93C2" ;
        when x"692" => cos_16 <= x"93A7" ;
        when x"693" => cos_16 <= x"938C" ;
        when x"694" => cos_16 <= x"9372" ;
        when x"695" => cos_16 <= x"9357" ;
        when x"696" => cos_16 <= x"933D" ;
        when x"697" => cos_16 <= x"9322" ;
        when x"698" => cos_16 <= x"9308" ;
        when x"699" => cos_16 <= x"92ED" ;
        when x"69A" => cos_16 <= x"92D3" ;
        when x"69B" => cos_16 <= x"92B9" ;
        when x"69C" => cos_16 <= x"929F" ;
        when x"69D" => cos_16 <= x"9285" ;
        when x"69E" => cos_16 <= x"926B" ;
        when x"69F" => cos_16 <= x"9251" ;
        when x"6A0" => cos_16 <= x"9237" ;
        when x"6A1" => cos_16 <= x"921D" ;
        when x"6A2" => cos_16 <= x"9203" ;
        when x"6A3" => cos_16 <= x"91EA" ;
        when x"6A4" => cos_16 <= x"91D0" ;
        when x"6A5" => cos_16 <= x"91B6" ;
        when x"6A6" => cos_16 <= x"919D" ;
        when x"6A7" => cos_16 <= x"9184" ;
        when x"6A8" => cos_16 <= x"916A" ;
        when x"6A9" => cos_16 <= x"9151" ;
        when x"6AA" => cos_16 <= x"9138" ;
        when x"6AB" => cos_16 <= x"911F" ;
        when x"6AC" => cos_16 <= x"9105" ;
        when x"6AD" => cos_16 <= x"90EC" ;
        when x"6AE" => cos_16 <= x"90D4" ;
        when x"6AF" => cos_16 <= x"90BB" ;
        when x"6B0" => cos_16 <= x"90A2" ;
        when x"6B1" => cos_16 <= x"9089" ;
        when x"6B2" => cos_16 <= x"9070" ;
        when x"6B3" => cos_16 <= x"9058" ;
        when x"6B4" => cos_16 <= x"903F" ;
        when x"6B5" => cos_16 <= x"9027" ;
        when x"6B6" => cos_16 <= x"900E" ;
        when x"6B7" => cos_16 <= x"8FF6" ;
        when x"6B8" => cos_16 <= x"8FDE" ;
        when x"6B9" => cos_16 <= x"8FC6" ;
        when x"6BA" => cos_16 <= x"8FAD" ;
        when x"6BB" => cos_16 <= x"8F95" ;
        when x"6BC" => cos_16 <= x"8F7D" ;
        when x"6BD" => cos_16 <= x"8F65" ;
        when x"6BE" => cos_16 <= x"8F4E" ;
        when x"6BF" => cos_16 <= x"8F36" ;
        when x"6C0" => cos_16 <= x"8F1E" ;
        when x"6C1" => cos_16 <= x"8F06" ;
        when x"6C2" => cos_16 <= x"8EEF" ;
        when x"6C3" => cos_16 <= x"8ED7" ;
        when x"6C4" => cos_16 <= x"8EC0" ;
        when x"6C5" => cos_16 <= x"8EA8" ;
        when x"6C6" => cos_16 <= x"8E91" ;
        when x"6C7" => cos_16 <= x"8E7A" ;
        when x"6C8" => cos_16 <= x"8E63" ;
        when x"6C9" => cos_16 <= x"8E4C" ;
        when x"6CA" => cos_16 <= x"8E35" ;
        when x"6CB" => cos_16 <= x"8E1E" ;
        when x"6CC" => cos_16 <= x"8E07" ;
        when x"6CD" => cos_16 <= x"8DF0" ;
        when x"6CE" => cos_16 <= x"8DD9" ;
        when x"6CF" => cos_16 <= x"8DC2" ;
        when x"6D0" => cos_16 <= x"8DAC" ;
        when x"6D1" => cos_16 <= x"8D95" ;
        when x"6D2" => cos_16 <= x"8D7F" ;
        when x"6D3" => cos_16 <= x"8D68" ;
        when x"6D4" => cos_16 <= x"8D52" ;
        when x"6D5" => cos_16 <= x"8D3C" ;
        when x"6D6" => cos_16 <= x"8D25" ;
        when x"6D7" => cos_16 <= x"8D0F" ;
        when x"6D8" => cos_16 <= x"8CF9" ;
        when x"6D9" => cos_16 <= x"8CE3" ;
        when x"6DA" => cos_16 <= x"8CCD" ;
        when x"6DB" => cos_16 <= x"8CB7" ;
        when x"6DC" => cos_16 <= x"8CA2" ;
        when x"6DD" => cos_16 <= x"8C8C" ;
        when x"6DE" => cos_16 <= x"8C76" ;
        when x"6DF" => cos_16 <= x"8C61" ;
        when x"6E0" => cos_16 <= x"8C4B" ;
        when x"6E1" => cos_16 <= x"8C36" ;
        when x"6E2" => cos_16 <= x"8C20" ;
        when x"6E3" => cos_16 <= x"8C0B" ;
        when x"6E4" => cos_16 <= x"8BF6" ;
        when x"6E5" => cos_16 <= x"8BE0" ;
        when x"6E6" => cos_16 <= x"8BCB" ;
        when x"6E7" => cos_16 <= x"8BB6" ;
        when x"6E8" => cos_16 <= x"8BA1" ;
        when x"6E9" => cos_16 <= x"8B8C" ;
        when x"6EA" => cos_16 <= x"8B78" ;
        when x"6EB" => cos_16 <= x"8B63" ;
        when x"6EC" => cos_16 <= x"8B4E" ;
        when x"6ED" => cos_16 <= x"8B3A" ;
        when x"6EE" => cos_16 <= x"8B25" ;
        when x"6EF" => cos_16 <= x"8B10" ;
        when x"6F0" => cos_16 <= x"8AFC" ;
        when x"6F1" => cos_16 <= x"8AE8" ;
        when x"6F2" => cos_16 <= x"8AD3" ;
        when x"6F3" => cos_16 <= x"8ABF" ;
        when x"6F4" => cos_16 <= x"8AAB" ;
        when x"6F5" => cos_16 <= x"8A97" ;
        when x"6F6" => cos_16 <= x"8A83" ;
        when x"6F7" => cos_16 <= x"8A6F" ;
        when x"6F8" => cos_16 <= x"8A5B" ;
        when x"6F9" => cos_16 <= x"8A48" ;
        when x"6FA" => cos_16 <= x"8A34" ;
        when x"6FB" => cos_16 <= x"8A20" ;
        when x"6FC" => cos_16 <= x"8A0D" ;
        when x"6FD" => cos_16 <= x"89F9" ;
        when x"6FE" => cos_16 <= x"89E6" ;
        when x"6FF" => cos_16 <= x"89D3" ;
        when x"700" => cos_16 <= x"89BF" ;
        when x"701" => cos_16 <= x"89AC" ;
        when x"702" => cos_16 <= x"8999" ;
        when x"703" => cos_16 <= x"8986" ;
        when x"704" => cos_16 <= x"8973" ;
        when x"705" => cos_16 <= x"8960" ;
        when x"706" => cos_16 <= x"894D" ;
        when x"707" => cos_16 <= x"893A" ;
        when x"708" => cos_16 <= x"8928" ;
        when x"709" => cos_16 <= x"8915" ;
        when x"70A" => cos_16 <= x"8902" ;
        when x"70B" => cos_16 <= x"88F0" ;
        when x"70C" => cos_16 <= x"88DE" ;
        when x"70D" => cos_16 <= x"88CB" ;
        when x"70E" => cos_16 <= x"88B9" ;
        when x"70F" => cos_16 <= x"88A7" ;
        when x"710" => cos_16 <= x"8895" ;
        when x"711" => cos_16 <= x"8883" ;
        when x"712" => cos_16 <= x"8871" ;
        when x"713" => cos_16 <= x"885F" ;
        when x"714" => cos_16 <= x"884D" ;
        when x"715" => cos_16 <= x"883B" ;
        when x"716" => cos_16 <= x"8829" ;
        when x"717" => cos_16 <= x"8818" ;
        when x"718" => cos_16 <= x"8806" ;
        when x"719" => cos_16 <= x"87F5" ;
        when x"71A" => cos_16 <= x"87E3" ;
        when x"71B" => cos_16 <= x"87D2" ;
        when x"71C" => cos_16 <= x"87C1" ;
        when x"71D" => cos_16 <= x"87B0" ;
        when x"71E" => cos_16 <= x"879E" ;
        when x"71F" => cos_16 <= x"878D" ;
        when x"720" => cos_16 <= x"877C" ;
        when x"721" => cos_16 <= x"876C" ;
        when x"722" => cos_16 <= x"875B" ;
        when x"723" => cos_16 <= x"874A" ;
        when x"724" => cos_16 <= x"8739" ;
        when x"725" => cos_16 <= x"8729" ;
        when x"726" => cos_16 <= x"8718" ;
        when x"727" => cos_16 <= x"8708" ;
        when x"728" => cos_16 <= x"86F7" ;
        when x"729" => cos_16 <= x"86E7" ;
        when x"72A" => cos_16 <= x"86D7" ;
        when x"72B" => cos_16 <= x"86C7" ;
        when x"72C" => cos_16 <= x"86B6" ;
        when x"72D" => cos_16 <= x"86A6" ;
        when x"72E" => cos_16 <= x"8696" ;
        when x"72F" => cos_16 <= x"8687" ;
        when x"730" => cos_16 <= x"8677" ;
        when x"731" => cos_16 <= x"8667" ;
        when x"732" => cos_16 <= x"8657" ;
        when x"733" => cos_16 <= x"8648" ;
        when x"734" => cos_16 <= x"8638" ;
        when x"735" => cos_16 <= x"8629" ;
        when x"736" => cos_16 <= x"861A" ;
        when x"737" => cos_16 <= x"860A" ;
        when x"738" => cos_16 <= x"85FB" ;
        when x"739" => cos_16 <= x"85EC" ;
        when x"73A" => cos_16 <= x"85DD" ;
        when x"73B" => cos_16 <= x"85CE" ;
        when x"73C" => cos_16 <= x"85BF" ;
        when x"73D" => cos_16 <= x"85B0" ;
        when x"73E" => cos_16 <= x"85A1" ;
        when x"73F" => cos_16 <= x"8593" ;
        when x"740" => cos_16 <= x"8584" ;
        when x"741" => cos_16 <= x"8575" ;
        when x"742" => cos_16 <= x"8567" ;
        when x"743" => cos_16 <= x"8558" ;
        when x"744" => cos_16 <= x"854A" ;
        when x"745" => cos_16 <= x"853C" ;
        when x"746" => cos_16 <= x"852E" ;
        when x"747" => cos_16 <= x"8520" ;
        when x"748" => cos_16 <= x"8512" ;
        when x"749" => cos_16 <= x"8504" ;
        when x"74A" => cos_16 <= x"84F6" ;
        when x"74B" => cos_16 <= x"84E8" ;
        when x"74C" => cos_16 <= x"84DA" ;
        when x"74D" => cos_16 <= x"84CD" ;
        when x"74E" => cos_16 <= x"84BF" ;
        when x"74F" => cos_16 <= x"84B1" ;
        when x"750" => cos_16 <= x"84A4" ;
        when x"751" => cos_16 <= x"8497" ;
        when x"752" => cos_16 <= x"8489" ;
        when x"753" => cos_16 <= x"847C" ;
        when x"754" => cos_16 <= x"846F" ;
        when x"755" => cos_16 <= x"8462" ;
        when x"756" => cos_16 <= x"8455" ;
        when x"757" => cos_16 <= x"8448" ;
        when x"758" => cos_16 <= x"843B" ;
        when x"759" => cos_16 <= x"842E" ;
        when x"75A" => cos_16 <= x"8422" ;
        when x"75B" => cos_16 <= x"8415" ;
        when x"75C" => cos_16 <= x"8408" ;
        when x"75D" => cos_16 <= x"83FC" ;
        when x"75E" => cos_16 <= x"83F0" ;
        when x"75F" => cos_16 <= x"83E3" ;
        when x"760" => cos_16 <= x"83D7" ;
        when x"761" => cos_16 <= x"83CB" ;
        when x"762" => cos_16 <= x"83BF" ;
        when x"763" => cos_16 <= x"83B3" ;
        when x"764" => cos_16 <= x"83A7" ;
        when x"765" => cos_16 <= x"839B" ;
        when x"766" => cos_16 <= x"838F" ;
        when x"767" => cos_16 <= x"8383" ;
        when x"768" => cos_16 <= x"8378" ;
        when x"769" => cos_16 <= x"836C" ;
        when x"76A" => cos_16 <= x"8361" ;
        when x"76B" => cos_16 <= x"8355" ;
        when x"76C" => cos_16 <= x"834A" ;
        when x"76D" => cos_16 <= x"833F" ;
        when x"76E" => cos_16 <= x"8333" ;
        when x"76F" => cos_16 <= x"8328" ;
        when x"770" => cos_16 <= x"831D" ;
        when x"771" => cos_16 <= x"8312" ;
        when x"772" => cos_16 <= x"8307" ;
        when x"773" => cos_16 <= x"82FC" ;
        when x"774" => cos_16 <= x"82F2" ;
        when x"775" => cos_16 <= x"82E7" ;
        when x"776" => cos_16 <= x"82DC" ;
        when x"777" => cos_16 <= x"82D2" ;
        when x"778" => cos_16 <= x"82C7" ;
        when x"779" => cos_16 <= x"82BD" ;
        when x"77A" => cos_16 <= x"82B3" ;
        when x"77B" => cos_16 <= x"82A9" ;
        when x"77C" => cos_16 <= x"829E" ;
        when x"77D" => cos_16 <= x"8294" ;
        when x"77E" => cos_16 <= x"828A" ;
        when x"77F" => cos_16 <= x"8280" ;
        when x"780" => cos_16 <= x"8277" ;
        when x"781" => cos_16 <= x"826D" ;
        when x"782" => cos_16 <= x"8263" ;
        when x"783" => cos_16 <= x"825A" ;
        when x"784" => cos_16 <= x"8250" ;
        when x"785" => cos_16 <= x"8247" ;
        when x"786" => cos_16 <= x"823D" ;
        when x"787" => cos_16 <= x"8234" ;
        when x"788" => cos_16 <= x"822B" ;
        when x"789" => cos_16 <= x"8221" ;
        when x"78A" => cos_16 <= x"8218" ;
        when x"78B" => cos_16 <= x"820F" ;
        when x"78C" => cos_16 <= x"8206" ;
        when x"78D" => cos_16 <= x"81FE" ;
        when x"78E" => cos_16 <= x"81F5" ;
        when x"78F" => cos_16 <= x"81EC" ;
        when x"790" => cos_16 <= x"81E3" ;
        when x"791" => cos_16 <= x"81DB" ;
        when x"792" => cos_16 <= x"81D2" ;
        when x"793" => cos_16 <= x"81CA" ;
        when x"794" => cos_16 <= x"81C2" ;
        when x"795" => cos_16 <= x"81B9" ;
        when x"796" => cos_16 <= x"81B1" ;
        when x"797" => cos_16 <= x"81A9" ;
        when x"798" => cos_16 <= x"81A1" ;
        when x"799" => cos_16 <= x"8199" ;
        when x"79A" => cos_16 <= x"8191" ;
        when x"79B" => cos_16 <= x"8189" ;
        when x"79C" => cos_16 <= x"8182" ;
        when x"79D" => cos_16 <= x"817A" ;
        when x"79E" => cos_16 <= x"8173" ;
        when x"79F" => cos_16 <= x"816B" ;
        when x"7A0" => cos_16 <= x"8164" ;
        when x"7A1" => cos_16 <= x"815C" ;
        when x"7A2" => cos_16 <= x"8155" ;
        when x"7A3" => cos_16 <= x"814E" ;
        when x"7A4" => cos_16 <= x"8147" ;
        when x"7A5" => cos_16 <= x"8140" ;
        when x"7A6" => cos_16 <= x"8139" ;
        when x"7A7" => cos_16 <= x"8132" ;
        when x"7A8" => cos_16 <= x"812B" ;
        when x"7A9" => cos_16 <= x"8124" ;
        when x"7AA" => cos_16 <= x"811E" ;
        when x"7AB" => cos_16 <= x"8117" ;
        when x"7AC" => cos_16 <= x"8111" ;
        when x"7AD" => cos_16 <= x"810A" ;
        when x"7AE" => cos_16 <= x"8104" ;
        when x"7AF" => cos_16 <= x"80FE" ;
        when x"7B0" => cos_16 <= x"80F7" ;
        when x"7B1" => cos_16 <= x"80F1" ;
        when x"7B2" => cos_16 <= x"80EB" ;
        when x"7B3" => cos_16 <= x"80E5" ;
        when x"7B4" => cos_16 <= x"80DF" ;
        when x"7B5" => cos_16 <= x"80DA" ;
        when x"7B6" => cos_16 <= x"80D4" ;
        when x"7B7" => cos_16 <= x"80CE" ;
        when x"7B8" => cos_16 <= x"80C9" ;
        when x"7B9" => cos_16 <= x"80C3" ;
        when x"7BA" => cos_16 <= x"80BE" ;
        when x"7BB" => cos_16 <= x"80B8" ;
        when x"7BC" => cos_16 <= x"80B3" ;
        when x"7BD" => cos_16 <= x"80AE" ;
        when x"7BE" => cos_16 <= x"80A9" ;
        when x"7BF" => cos_16 <= x"80A4" ;
        when x"7C0" => cos_16 <= x"809F" ;
        when x"7C1" => cos_16 <= x"809A" ;
        when x"7C2" => cos_16 <= x"8095" ;
        when x"7C3" => cos_16 <= x"8090" ;
        when x"7C4" => cos_16 <= x"808C" ;
        when x"7C5" => cos_16 <= x"8087" ;
        when x"7C6" => cos_16 <= x"8083" ;
        when x"7C7" => cos_16 <= x"807E" ;
        when x"7C8" => cos_16 <= x"807A" ;
        when x"7C9" => cos_16 <= x"8076" ;
        when x"7CA" => cos_16 <= x"8071" ;
        when x"7CB" => cos_16 <= x"806D" ;
        when x"7CC" => cos_16 <= x"8069" ;
        when x"7CD" => cos_16 <= x"8065" ;
        when x"7CE" => cos_16 <= x"8061" ;
        when x"7CF" => cos_16 <= x"805E" ;
        when x"7D0" => cos_16 <= x"805A" ;
        when x"7D1" => cos_16 <= x"8056" ;
        when x"7D2" => cos_16 <= x"8053" ;
        when x"7D3" => cos_16 <= x"804F" ;
        when x"7D4" => cos_16 <= x"804C" ;
        when x"7D5" => cos_16 <= x"8048" ;
        when x"7D6" => cos_16 <= x"8045" ;
        when x"7D7" => cos_16 <= x"8042" ;
        when x"7D8" => cos_16 <= x"803F" ;
        when x"7D9" => cos_16 <= x"803C" ;
        when x"7DA" => cos_16 <= x"8039" ;
        when x"7DB" => cos_16 <= x"8036" ;
        when x"7DC" => cos_16 <= x"8033" ;
        when x"7DD" => cos_16 <= x"8030" ;
        when x"7DE" => cos_16 <= x"802E" ;
        when x"7DF" => cos_16 <= x"802B" ;
        when x"7E0" => cos_16 <= x"8028" ;
        when x"7E1" => cos_16 <= x"8026" ;
        when x"7E2" => cos_16 <= x"8024" ;
        when x"7E3" => cos_16 <= x"8021" ;
        when x"7E4" => cos_16 <= x"801F" ;
        when x"7E5" => cos_16 <= x"801D" ;
        when x"7E6" => cos_16 <= x"801B" ;
        when x"7E7" => cos_16 <= x"8019" ;
        when x"7E8" => cos_16 <= x"8017" ;
        when x"7E9" => cos_16 <= x"8015" ;
        when x"7EA" => cos_16 <= x"8014" ;
        when x"7EB" => cos_16 <= x"8012" ;
        when x"7EC" => cos_16 <= x"8010" ;
        when x"7ED" => cos_16 <= x"800F" ;
        when x"7EE" => cos_16 <= x"800D" ;
        when x"7EF" => cos_16 <= x"800C" ;
        when x"7F0" => cos_16 <= x"800B" ;
        when x"7F1" => cos_16 <= x"800A" ;
        when x"7F2" => cos_16 <= x"8009" ;
        when x"7F3" => cos_16 <= x"8008" ;
        when x"7F4" => cos_16 <= x"8007" ;
        when x"7F5" => cos_16 <= x"8006" ;
        when x"7F6" => cos_16 <= x"8005" ;
        when x"7F7" => cos_16 <= x"8004" ;
        when x"7F8" => cos_16 <= x"8003" ;
        when x"7F9" => cos_16 <= x"8003" ;
        when x"7FA" => cos_16 <= x"8002" ;
        when x"7FB" => cos_16 <= x"8002" ;
        when x"7FC" => cos_16 <= x"8002" ;
        when x"7FD" => cos_16 <= x"8001" ;
        when x"7FE" => cos_16 <= x"8001" ;
        when x"7FF" => cos_16 <= x"8001" ;
        when x"800" => cos_16 <= x"8001" ;
        when x"801" => cos_16 <= x"8001" ;
        when x"802" => cos_16 <= x"8001" ;
        when x"803" => cos_16 <= x"8001" ;
        when x"804" => cos_16 <= x"8002" ;
        when x"805" => cos_16 <= x"8002" ;
        when x"806" => cos_16 <= x"8002" ;
        when x"807" => cos_16 <= x"8003" ;
        when x"808" => cos_16 <= x"8003" ;
        when x"809" => cos_16 <= x"8004" ;
        when x"80A" => cos_16 <= x"8005" ;
        when x"80B" => cos_16 <= x"8006" ;
        when x"80C" => cos_16 <= x"8007" ;
        when x"80D" => cos_16 <= x"8008" ;
        when x"80E" => cos_16 <= x"8009" ;
        when x"80F" => cos_16 <= x"800A" ;
        when x"810" => cos_16 <= x"800B" ;
        when x"811" => cos_16 <= x"800C" ;
        when x"812" => cos_16 <= x"800D" ;
        when x"813" => cos_16 <= x"800F" ;
        when x"814" => cos_16 <= x"8010" ;
        when x"815" => cos_16 <= x"8012" ;
        when x"816" => cos_16 <= x"8014" ;
        when x"817" => cos_16 <= x"8015" ;
        when x"818" => cos_16 <= x"8017" ;
        when x"819" => cos_16 <= x"8019" ;
        when x"81A" => cos_16 <= x"801B" ;
        when x"81B" => cos_16 <= x"801D" ;
        when x"81C" => cos_16 <= x"801F" ;
        when x"81D" => cos_16 <= x"8021" ;
        when x"81E" => cos_16 <= x"8024" ;
        when x"81F" => cos_16 <= x"8026" ;
        when x"820" => cos_16 <= x"8028" ;
        when x"821" => cos_16 <= x"802B" ;
        when x"822" => cos_16 <= x"802E" ;
        when x"823" => cos_16 <= x"8030" ;
        when x"824" => cos_16 <= x"8033" ;
        when x"825" => cos_16 <= x"8036" ;
        when x"826" => cos_16 <= x"8039" ;
        when x"827" => cos_16 <= x"803C" ;
        when x"828" => cos_16 <= x"803F" ;
        when x"829" => cos_16 <= x"8042" ;
        when x"82A" => cos_16 <= x"8045" ;
        when x"82B" => cos_16 <= x"8048" ;
        when x"82C" => cos_16 <= x"804C" ;
        when x"82D" => cos_16 <= x"804F" ;
        when x"82E" => cos_16 <= x"8053" ;
        when x"82F" => cos_16 <= x"8056" ;
        when x"830" => cos_16 <= x"805A" ;
        when x"831" => cos_16 <= x"805E" ;
        when x"832" => cos_16 <= x"8061" ;
        when x"833" => cos_16 <= x"8065" ;
        when x"834" => cos_16 <= x"8069" ;
        when x"835" => cos_16 <= x"806D" ;
        when x"836" => cos_16 <= x"8071" ;
        when x"837" => cos_16 <= x"8076" ;
        when x"838" => cos_16 <= x"807A" ;
        when x"839" => cos_16 <= x"807E" ;
        when x"83A" => cos_16 <= x"8083" ;
        when x"83B" => cos_16 <= x"8087" ;
        when x"83C" => cos_16 <= x"808C" ;
        when x"83D" => cos_16 <= x"8090" ;
        when x"83E" => cos_16 <= x"8095" ;
        when x"83F" => cos_16 <= x"809A" ;
        when x"840" => cos_16 <= x"809F" ;
        when x"841" => cos_16 <= x"80A4" ;
        when x"842" => cos_16 <= x"80A9" ;
        when x"843" => cos_16 <= x"80AE" ;
        when x"844" => cos_16 <= x"80B3" ;
        when x"845" => cos_16 <= x"80B8" ;
        when x"846" => cos_16 <= x"80BE" ;
        when x"847" => cos_16 <= x"80C3" ;
        when x"848" => cos_16 <= x"80C9" ;
        when x"849" => cos_16 <= x"80CE" ;
        when x"84A" => cos_16 <= x"80D4" ;
        when x"84B" => cos_16 <= x"80DA" ;
        when x"84C" => cos_16 <= x"80DF" ;
        when x"84D" => cos_16 <= x"80E5" ;
        when x"84E" => cos_16 <= x"80EB" ;
        when x"84F" => cos_16 <= x"80F1" ;
        when x"850" => cos_16 <= x"80F7" ;
        when x"851" => cos_16 <= x"80FE" ;
        when x"852" => cos_16 <= x"8104" ;
        when x"853" => cos_16 <= x"810A" ;
        when x"854" => cos_16 <= x"8111" ;
        when x"855" => cos_16 <= x"8117" ;
        when x"856" => cos_16 <= x"811E" ;
        when x"857" => cos_16 <= x"8124" ;
        when x"858" => cos_16 <= x"812B" ;
        when x"859" => cos_16 <= x"8132" ;
        when x"85A" => cos_16 <= x"8139" ;
        when x"85B" => cos_16 <= x"8140" ;
        when x"85C" => cos_16 <= x"8147" ;
        when x"85D" => cos_16 <= x"814E" ;
        when x"85E" => cos_16 <= x"8155" ;
        when x"85F" => cos_16 <= x"815C" ;
        when x"860" => cos_16 <= x"8164" ;
        when x"861" => cos_16 <= x"816B" ;
        when x"862" => cos_16 <= x"8173" ;
        when x"863" => cos_16 <= x"817A" ;
        when x"864" => cos_16 <= x"8182" ;
        when x"865" => cos_16 <= x"8189" ;
        when x"866" => cos_16 <= x"8191" ;
        when x"867" => cos_16 <= x"8199" ;
        when x"868" => cos_16 <= x"81A1" ;
        when x"869" => cos_16 <= x"81A9" ;
        when x"86A" => cos_16 <= x"81B1" ;
        when x"86B" => cos_16 <= x"81B9" ;
        when x"86C" => cos_16 <= x"81C2" ;
        when x"86D" => cos_16 <= x"81CA" ;
        when x"86E" => cos_16 <= x"81D2" ;
        when x"86F" => cos_16 <= x"81DB" ;
        when x"870" => cos_16 <= x"81E3" ;
        when x"871" => cos_16 <= x"81EC" ;
        when x"872" => cos_16 <= x"81F5" ;
        when x"873" => cos_16 <= x"81FE" ;
        when x"874" => cos_16 <= x"8206" ;
        when x"875" => cos_16 <= x"820F" ;
        when x"876" => cos_16 <= x"8218" ;
        when x"877" => cos_16 <= x"8221" ;
        when x"878" => cos_16 <= x"822B" ;
        when x"879" => cos_16 <= x"8234" ;
        when x"87A" => cos_16 <= x"823D" ;
        when x"87B" => cos_16 <= x"8247" ;
        when x"87C" => cos_16 <= x"8250" ;
        when x"87D" => cos_16 <= x"825A" ;
        when x"87E" => cos_16 <= x"8263" ;
        when x"87F" => cos_16 <= x"826D" ;
        when x"880" => cos_16 <= x"8277" ;
        when x"881" => cos_16 <= x"8280" ;
        when x"882" => cos_16 <= x"828A" ;
        when x"883" => cos_16 <= x"8294" ;
        when x"884" => cos_16 <= x"829E" ;
        when x"885" => cos_16 <= x"82A9" ;
        when x"886" => cos_16 <= x"82B3" ;
        when x"887" => cos_16 <= x"82BD" ;
        when x"888" => cos_16 <= x"82C7" ;
        when x"889" => cos_16 <= x"82D2" ;
        when x"88A" => cos_16 <= x"82DC" ;
        when x"88B" => cos_16 <= x"82E7" ;
        when x"88C" => cos_16 <= x"82F2" ;
        when x"88D" => cos_16 <= x"82FC" ;
        when x"88E" => cos_16 <= x"8307" ;
        when x"88F" => cos_16 <= x"8312" ;
        when x"890" => cos_16 <= x"831D" ;
        when x"891" => cos_16 <= x"8328" ;
        when x"892" => cos_16 <= x"8333" ;
        when x"893" => cos_16 <= x"833F" ;
        when x"894" => cos_16 <= x"834A" ;
        when x"895" => cos_16 <= x"8355" ;
        when x"896" => cos_16 <= x"8361" ;
        when x"897" => cos_16 <= x"836C" ;
        when x"898" => cos_16 <= x"8378" ;
        when x"899" => cos_16 <= x"8383" ;
        when x"89A" => cos_16 <= x"838F" ;
        when x"89B" => cos_16 <= x"839B" ;
        when x"89C" => cos_16 <= x"83A7" ;
        when x"89D" => cos_16 <= x"83B3" ;
        when x"89E" => cos_16 <= x"83BF" ;
        when x"89F" => cos_16 <= x"83CB" ;
        when x"8A0" => cos_16 <= x"83D7" ;
        when x"8A1" => cos_16 <= x"83E3" ;
        when x"8A2" => cos_16 <= x"83F0" ;
        when x"8A3" => cos_16 <= x"83FC" ;
        when x"8A4" => cos_16 <= x"8408" ;
        when x"8A5" => cos_16 <= x"8415" ;
        when x"8A6" => cos_16 <= x"8422" ;
        when x"8A7" => cos_16 <= x"842E" ;
        when x"8A8" => cos_16 <= x"843B" ;
        when x"8A9" => cos_16 <= x"8448" ;
        when x"8AA" => cos_16 <= x"8455" ;
        when x"8AB" => cos_16 <= x"8462" ;
        when x"8AC" => cos_16 <= x"846F" ;
        when x"8AD" => cos_16 <= x"847C" ;
        when x"8AE" => cos_16 <= x"8489" ;
        when x"8AF" => cos_16 <= x"8497" ;
        when x"8B0" => cos_16 <= x"84A4" ;
        when x"8B1" => cos_16 <= x"84B1" ;
        when x"8B2" => cos_16 <= x"84BF" ;
        when x"8B3" => cos_16 <= x"84CD" ;
        when x"8B4" => cos_16 <= x"84DA" ;
        when x"8B5" => cos_16 <= x"84E8" ;
        when x"8B6" => cos_16 <= x"84F6" ;
        when x"8B7" => cos_16 <= x"8504" ;
        when x"8B8" => cos_16 <= x"8512" ;
        when x"8B9" => cos_16 <= x"8520" ;
        when x"8BA" => cos_16 <= x"852E" ;
        when x"8BB" => cos_16 <= x"853C" ;
        when x"8BC" => cos_16 <= x"854A" ;
        when x"8BD" => cos_16 <= x"8558" ;
        when x"8BE" => cos_16 <= x"8567" ;
        when x"8BF" => cos_16 <= x"8575" ;
        when x"8C0" => cos_16 <= x"8584" ;
        when x"8C1" => cos_16 <= x"8593" ;
        when x"8C2" => cos_16 <= x"85A1" ;
        when x"8C3" => cos_16 <= x"85B0" ;
        when x"8C4" => cos_16 <= x"85BF" ;
        when x"8C5" => cos_16 <= x"85CE" ;
        when x"8C6" => cos_16 <= x"85DD" ;
        when x"8C7" => cos_16 <= x"85EC" ;
        when x"8C8" => cos_16 <= x"85FB" ;
        when x"8C9" => cos_16 <= x"860A" ;
        when x"8CA" => cos_16 <= x"861A" ;
        when x"8CB" => cos_16 <= x"8629" ;
        when x"8CC" => cos_16 <= x"8638" ;
        when x"8CD" => cos_16 <= x"8648" ;
        when x"8CE" => cos_16 <= x"8657" ;
        when x"8CF" => cos_16 <= x"8667" ;
        when x"8D0" => cos_16 <= x"8677" ;
        when x"8D1" => cos_16 <= x"8687" ;
        when x"8D2" => cos_16 <= x"8696" ;
        when x"8D3" => cos_16 <= x"86A6" ;
        when x"8D4" => cos_16 <= x"86B6" ;
        when x"8D5" => cos_16 <= x"86C7" ;
        when x"8D6" => cos_16 <= x"86D7" ;
        when x"8D7" => cos_16 <= x"86E7" ;
        when x"8D8" => cos_16 <= x"86F7" ;
        when x"8D9" => cos_16 <= x"8708" ;
        when x"8DA" => cos_16 <= x"8718" ;
        when x"8DB" => cos_16 <= x"8729" ;
        when x"8DC" => cos_16 <= x"8739" ;
        when x"8DD" => cos_16 <= x"874A" ;
        when x"8DE" => cos_16 <= x"875B" ;
        when x"8DF" => cos_16 <= x"876C" ;
        when x"8E0" => cos_16 <= x"877C" ;
        when x"8E1" => cos_16 <= x"878D" ;
        when x"8E2" => cos_16 <= x"879E" ;
        when x"8E3" => cos_16 <= x"87B0" ;
        when x"8E4" => cos_16 <= x"87C1" ;
        when x"8E5" => cos_16 <= x"87D2" ;
        when x"8E6" => cos_16 <= x"87E3" ;
        when x"8E7" => cos_16 <= x"87F5" ;
        when x"8E8" => cos_16 <= x"8806" ;
        when x"8E9" => cos_16 <= x"8818" ;
        when x"8EA" => cos_16 <= x"8829" ;
        when x"8EB" => cos_16 <= x"883B" ;
        when x"8EC" => cos_16 <= x"884D" ;
        when x"8ED" => cos_16 <= x"885F" ;
        when x"8EE" => cos_16 <= x"8871" ;
        when x"8EF" => cos_16 <= x"8883" ;
        when x"8F0" => cos_16 <= x"8895" ;
        when x"8F1" => cos_16 <= x"88A7" ;
        when x"8F2" => cos_16 <= x"88B9" ;
        when x"8F3" => cos_16 <= x"88CB" ;
        when x"8F4" => cos_16 <= x"88DE" ;
        when x"8F5" => cos_16 <= x"88F0" ;
        when x"8F6" => cos_16 <= x"8902" ;
        when x"8F7" => cos_16 <= x"8915" ;
        when x"8F8" => cos_16 <= x"8928" ;
        when x"8F9" => cos_16 <= x"893A" ;
        when x"8FA" => cos_16 <= x"894D" ;
        when x"8FB" => cos_16 <= x"8960" ;
        when x"8FC" => cos_16 <= x"8973" ;
        when x"8FD" => cos_16 <= x"8986" ;
        when x"8FE" => cos_16 <= x"8999" ;
        when x"8FF" => cos_16 <= x"89AC" ;
        when x"900" => cos_16 <= x"89BF" ;
        when x"901" => cos_16 <= x"89D3" ;
        when x"902" => cos_16 <= x"89E6" ;
        when x"903" => cos_16 <= x"89F9" ;
        when x"904" => cos_16 <= x"8A0D" ;
        when x"905" => cos_16 <= x"8A20" ;
        when x"906" => cos_16 <= x"8A34" ;
        when x"907" => cos_16 <= x"8A48" ;
        when x"908" => cos_16 <= x"8A5B" ;
        when x"909" => cos_16 <= x"8A6F" ;
        when x"90A" => cos_16 <= x"8A83" ;
        when x"90B" => cos_16 <= x"8A97" ;
        when x"90C" => cos_16 <= x"8AAB" ;
        when x"90D" => cos_16 <= x"8ABF" ;
        when x"90E" => cos_16 <= x"8AD3" ;
        when x"90F" => cos_16 <= x"8AE8" ;
        when x"910" => cos_16 <= x"8AFC" ;
        when x"911" => cos_16 <= x"8B10" ;
        when x"912" => cos_16 <= x"8B25" ;
        when x"913" => cos_16 <= x"8B3A" ;
        when x"914" => cos_16 <= x"8B4E" ;
        when x"915" => cos_16 <= x"8B63" ;
        when x"916" => cos_16 <= x"8B78" ;
        when x"917" => cos_16 <= x"8B8C" ;
        when x"918" => cos_16 <= x"8BA1" ;
        when x"919" => cos_16 <= x"8BB6" ;
        when x"91A" => cos_16 <= x"8BCB" ;
        when x"91B" => cos_16 <= x"8BE0" ;
        when x"91C" => cos_16 <= x"8BF6" ;
        when x"91D" => cos_16 <= x"8C0B" ;
        when x"91E" => cos_16 <= x"8C20" ;
        when x"91F" => cos_16 <= x"8C36" ;
        when x"920" => cos_16 <= x"8C4B" ;
        when x"921" => cos_16 <= x"8C61" ;
        when x"922" => cos_16 <= x"8C76" ;
        when x"923" => cos_16 <= x"8C8C" ;
        when x"924" => cos_16 <= x"8CA2" ;
        when x"925" => cos_16 <= x"8CB7" ;
        when x"926" => cos_16 <= x"8CCD" ;
        when x"927" => cos_16 <= x"8CE3" ;
        when x"928" => cos_16 <= x"8CF9" ;
        when x"929" => cos_16 <= x"8D0F" ;
        when x"92A" => cos_16 <= x"8D25" ;
        when x"92B" => cos_16 <= x"8D3C" ;
        when x"92C" => cos_16 <= x"8D52" ;
        when x"92D" => cos_16 <= x"8D68" ;
        when x"92E" => cos_16 <= x"8D7F" ;
        when x"92F" => cos_16 <= x"8D95" ;
        when x"930" => cos_16 <= x"8DAC" ;
        when x"931" => cos_16 <= x"8DC2" ;
        when x"932" => cos_16 <= x"8DD9" ;
        when x"933" => cos_16 <= x"8DF0" ;
        when x"934" => cos_16 <= x"8E07" ;
        when x"935" => cos_16 <= x"8E1E" ;
        when x"936" => cos_16 <= x"8E35" ;
        when x"937" => cos_16 <= x"8E4C" ;
        when x"938" => cos_16 <= x"8E63" ;
        when x"939" => cos_16 <= x"8E7A" ;
        when x"93A" => cos_16 <= x"8E91" ;
        when x"93B" => cos_16 <= x"8EA8" ;
        when x"93C" => cos_16 <= x"8EC0" ;
        when x"93D" => cos_16 <= x"8ED7" ;
        when x"93E" => cos_16 <= x"8EEF" ;
        when x"93F" => cos_16 <= x"8F06" ;
        when x"940" => cos_16 <= x"8F1E" ;
        when x"941" => cos_16 <= x"8F36" ;
        when x"942" => cos_16 <= x"8F4E" ;
        when x"943" => cos_16 <= x"8F65" ;
        when x"944" => cos_16 <= x"8F7D" ;
        when x"945" => cos_16 <= x"8F95" ;
        when x"946" => cos_16 <= x"8FAD" ;
        when x"947" => cos_16 <= x"8FC6" ;
        when x"948" => cos_16 <= x"8FDE" ;
        when x"949" => cos_16 <= x"8FF6" ;
        when x"94A" => cos_16 <= x"900E" ;
        when x"94B" => cos_16 <= x"9027" ;
        when x"94C" => cos_16 <= x"903F" ;
        when x"94D" => cos_16 <= x"9058" ;
        when x"94E" => cos_16 <= x"9070" ;
        when x"94F" => cos_16 <= x"9089" ;
        when x"950" => cos_16 <= x"90A2" ;
        when x"951" => cos_16 <= x"90BB" ;
        when x"952" => cos_16 <= x"90D4" ;
        when x"953" => cos_16 <= x"90EC" ;
        when x"954" => cos_16 <= x"9105" ;
        when x"955" => cos_16 <= x"911F" ;
        when x"956" => cos_16 <= x"9138" ;
        when x"957" => cos_16 <= x"9151" ;
        when x"958" => cos_16 <= x"916A" ;
        when x"959" => cos_16 <= x"9184" ;
        when x"95A" => cos_16 <= x"919D" ;
        when x"95B" => cos_16 <= x"91B6" ;
        when x"95C" => cos_16 <= x"91D0" ;
        when x"95D" => cos_16 <= x"91EA" ;
        when x"95E" => cos_16 <= x"9203" ;
        when x"95F" => cos_16 <= x"921D" ;
        when x"960" => cos_16 <= x"9237" ;
        when x"961" => cos_16 <= x"9251" ;
        when x"962" => cos_16 <= x"926B" ;
        when x"963" => cos_16 <= x"9285" ;
        when x"964" => cos_16 <= x"929F" ;
        when x"965" => cos_16 <= x"92B9" ;
        when x"966" => cos_16 <= x"92D3" ;
        when x"967" => cos_16 <= x"92ED" ;
        when x"968" => cos_16 <= x"9308" ;
        when x"969" => cos_16 <= x"9322" ;
        when x"96A" => cos_16 <= x"933D" ;
        when x"96B" => cos_16 <= x"9357" ;
        when x"96C" => cos_16 <= x"9372" ;
        when x"96D" => cos_16 <= x"938C" ;
        when x"96E" => cos_16 <= x"93A7" ;
        when x"96F" => cos_16 <= x"93C2" ;
        when x"970" => cos_16 <= x"93DD" ;
        when x"971" => cos_16 <= x"93F8" ;
        when x"972" => cos_16 <= x"9413" ;
        when x"973" => cos_16 <= x"942E" ;
        when x"974" => cos_16 <= x"9449" ;
        when x"975" => cos_16 <= x"9464" ;
        when x"976" => cos_16 <= x"947F" ;
        when x"977" => cos_16 <= x"949B" ;
        when x"978" => cos_16 <= x"94B6" ;
        when x"979" => cos_16 <= x"94D1" ;
        when x"97A" => cos_16 <= x"94ED" ;
        when x"97B" => cos_16 <= x"9508" ;
        when x"97C" => cos_16 <= x"9524" ;
        when x"97D" => cos_16 <= x"9540" ;
        when x"97E" => cos_16 <= x"955C" ;
        when x"97F" => cos_16 <= x"9577" ;
        when x"980" => cos_16 <= x"9593" ;
        when x"981" => cos_16 <= x"95AF" ;
        when x"982" => cos_16 <= x"95CB" ;
        when x"983" => cos_16 <= x"95E7" ;
        when x"984" => cos_16 <= x"9603" ;
        when x"985" => cos_16 <= x"9620" ;
        when x"986" => cos_16 <= x"963C" ;
        when x"987" => cos_16 <= x"9658" ;
        when x"988" => cos_16 <= x"9675" ;
        when x"989" => cos_16 <= x"9691" ;
        when x"98A" => cos_16 <= x"96AE" ;
        when x"98B" => cos_16 <= x"96CA" ;
        when x"98C" => cos_16 <= x"96E7" ;
        when x"98D" => cos_16 <= x"9704" ;
        when x"98E" => cos_16 <= x"9720" ;
        when x"98F" => cos_16 <= x"973D" ;
        when x"990" => cos_16 <= x"975A" ;
        when x"991" => cos_16 <= x"9777" ;
        when x"992" => cos_16 <= x"9794" ;
        when x"993" => cos_16 <= x"97B1" ;
        when x"994" => cos_16 <= x"97CE" ;
        when x"995" => cos_16 <= x"97EC" ;
        when x"996" => cos_16 <= x"9809" ;
        when x"997" => cos_16 <= x"9826" ;
        when x"998" => cos_16 <= x"9844" ;
        when x"999" => cos_16 <= x"9861" ;
        when x"99A" => cos_16 <= x"987F" ;
        when x"99B" => cos_16 <= x"989C" ;
        when x"99C" => cos_16 <= x"98BA" ;
        when x"99D" => cos_16 <= x"98D8" ;
        when x"99E" => cos_16 <= x"98F6" ;
        when x"99F" => cos_16 <= x"9913" ;
        when x"9A0" => cos_16 <= x"9931" ;
        when x"9A1" => cos_16 <= x"994F" ;
        when x"9A2" => cos_16 <= x"996D" ;
        when x"9A3" => cos_16 <= x"998B" ;
        when x"9A4" => cos_16 <= x"99AA" ;
        when x"9A5" => cos_16 <= x"99C8" ;
        when x"9A6" => cos_16 <= x"99E6" ;
        when x"9A7" => cos_16 <= x"9A04" ;
        when x"9A8" => cos_16 <= x"9A23" ;
        when x"9A9" => cos_16 <= x"9A41" ;
        when x"9AA" => cos_16 <= x"9A60" ;
        when x"9AB" => cos_16 <= x"9A7E" ;
        when x"9AC" => cos_16 <= x"9A9D" ;
        when x"9AD" => cos_16 <= x"9ABC" ;
        when x"9AE" => cos_16 <= x"9ADB" ;
        when x"9AF" => cos_16 <= x"9AF9" ;
        when x"9B0" => cos_16 <= x"9B18" ;
        when x"9B1" => cos_16 <= x"9B37" ;
        when x"9B2" => cos_16 <= x"9B56" ;
        when x"9B3" => cos_16 <= x"9B75" ;
        when x"9B4" => cos_16 <= x"9B94" ;
        when x"9B5" => cos_16 <= x"9BB4" ;
        when x"9B6" => cos_16 <= x"9BD3" ;
        when x"9B7" => cos_16 <= x"9BF2" ;
        when x"9B8" => cos_16 <= x"9C12" ;
        when x"9B9" => cos_16 <= x"9C31" ;
        when x"9BA" => cos_16 <= x"9C51" ;
        when x"9BB" => cos_16 <= x"9C70" ;
        when x"9BC" => cos_16 <= x"9C90" ;
        when x"9BD" => cos_16 <= x"9CAF" ;
        when x"9BE" => cos_16 <= x"9CCF" ;
        when x"9BF" => cos_16 <= x"9CEF" ;
        when x"9C0" => cos_16 <= x"9D0F" ;
        when x"9C1" => cos_16 <= x"9D2F" ;
        when x"9C2" => cos_16 <= x"9D4F" ;
        when x"9C3" => cos_16 <= x"9D6F" ;
        when x"9C4" => cos_16 <= x"9D8F" ;
        when x"9C5" => cos_16 <= x"9DAF" ;
        when x"9C6" => cos_16 <= x"9DCF" ;
        when x"9C7" => cos_16 <= x"9DEF" ;
        when x"9C8" => cos_16 <= x"9E10" ;
        when x"9C9" => cos_16 <= x"9E30" ;
        when x"9CA" => cos_16 <= x"9E51" ;
        when x"9CB" => cos_16 <= x"9E71" ;
        when x"9CC" => cos_16 <= x"9E92" ;
        when x"9CD" => cos_16 <= x"9EB2" ;
        when x"9CE" => cos_16 <= x"9ED3" ;
        when x"9CF" => cos_16 <= x"9EF4" ;
        when x"9D0" => cos_16 <= x"9F15" ;
        when x"9D1" => cos_16 <= x"9F35" ;
        when x"9D2" => cos_16 <= x"9F56" ;
        when x"9D3" => cos_16 <= x"9F77" ;
        when x"9D4" => cos_16 <= x"9F98" ;
        when x"9D5" => cos_16 <= x"9FB9" ;
        when x"9D6" => cos_16 <= x"9FDB" ;
        when x"9D7" => cos_16 <= x"9FFC" ;
        when x"9D8" => cos_16 <= x"A01D" ;
        when x"9D9" => cos_16 <= x"A03E" ;
        when x"9DA" => cos_16 <= x"A060" ;
        when x"9DB" => cos_16 <= x"A081" ;
        when x"9DC" => cos_16 <= x"A0A3" ;
        when x"9DD" => cos_16 <= x"A0C4" ;
        when x"9DE" => cos_16 <= x"A0E6" ;
        when x"9DF" => cos_16 <= x"A108" ;
        when x"9E0" => cos_16 <= x"A129" ;
        when x"9E1" => cos_16 <= x"A14B" ;
        when x"9E2" => cos_16 <= x"A16D" ;
        when x"9E3" => cos_16 <= x"A18F" ;
        when x"9E4" => cos_16 <= x"A1B1" ;
        when x"9E5" => cos_16 <= x"A1D3" ;
        when x"9E6" => cos_16 <= x"A1F5" ;
        when x"9E7" => cos_16 <= x"A217" ;
        when x"9E8" => cos_16 <= x"A239" ;
        when x"9E9" => cos_16 <= x"A25B" ;
        when x"9EA" => cos_16 <= x"A27E" ;
        when x"9EB" => cos_16 <= x"A2A0" ;
        when x"9EC" => cos_16 <= x"A2C2" ;
        when x"9ED" => cos_16 <= x"A2E5" ;
        when x"9EE" => cos_16 <= x"A307" ;
        when x"9EF" => cos_16 <= x"A32A" ;
        when x"9F0" => cos_16 <= x"A34D" ;
        when x"9F1" => cos_16 <= x"A36F" ;
        when x"9F2" => cos_16 <= x"A392" ;
        when x"9F3" => cos_16 <= x"A3B5" ;
        when x"9F4" => cos_16 <= x"A3D8" ;
        when x"9F5" => cos_16 <= x"A3FB" ;
        when x"9F6" => cos_16 <= x"A41E" ;
        when x"9F7" => cos_16 <= x"A441" ;
        when x"9F8" => cos_16 <= x"A464" ;
        when x"9F9" => cos_16 <= x"A487" ;
        when x"9FA" => cos_16 <= x"A4AA" ;
        when x"9FB" => cos_16 <= x"A4CD" ;
        when x"9FC" => cos_16 <= x"A4F1" ;
        when x"9FD" => cos_16 <= x"A514" ;
        when x"9FE" => cos_16 <= x"A537" ;
        when x"9FF" => cos_16 <= x"A55B" ;
        when x"A00" => cos_16 <= x"A57E" ;
        when x"A01" => cos_16 <= x"A5A2" ;
        when x"A02" => cos_16 <= x"A5C5" ;
        when x"A03" => cos_16 <= x"A5E9" ;
        when x"A04" => cos_16 <= x"A60D" ;
        when x"A05" => cos_16 <= x"A631" ;
        when x"A06" => cos_16 <= x"A654" ;
        when x"A07" => cos_16 <= x"A678" ;
        when x"A08" => cos_16 <= x"A69C" ;
        when x"A09" => cos_16 <= x"A6C0" ;
        when x"A0A" => cos_16 <= x"A6E4" ;
        when x"A0B" => cos_16 <= x"A708" ;
        when x"A0C" => cos_16 <= x"A72D" ;
        when x"A0D" => cos_16 <= x"A751" ;
        when x"A0E" => cos_16 <= x"A775" ;
        when x"A0F" => cos_16 <= x"A799" ;
        when x"A10" => cos_16 <= x"A7BE" ;
        when x"A11" => cos_16 <= x"A7E2" ;
        when x"A12" => cos_16 <= x"A807" ;
        when x"A13" => cos_16 <= x"A82B" ;
        when x"A14" => cos_16 <= x"A850" ;
        when x"A15" => cos_16 <= x"A875" ;
        when x"A16" => cos_16 <= x"A899" ;
        when x"A17" => cos_16 <= x"A8BE" ;
        when x"A18" => cos_16 <= x"A8E3" ;
        when x"A19" => cos_16 <= x"A908" ;
        when x"A1A" => cos_16 <= x"A92D" ;
        when x"A1B" => cos_16 <= x"A951" ;
        when x"A1C" => cos_16 <= x"A976" ;
        when x"A1D" => cos_16 <= x"A99C" ;
        when x"A1E" => cos_16 <= x"A9C1" ;
        when x"A1F" => cos_16 <= x"A9E6" ;
        when x"A20" => cos_16 <= x"AA0B" ;
        when x"A21" => cos_16 <= x"AA30" ;
        when x"A22" => cos_16 <= x"AA56" ;
        when x"A23" => cos_16 <= x"AA7B" ;
        when x"A24" => cos_16 <= x"AAA0" ;
        when x"A25" => cos_16 <= x"AAC6" ;
        when x"A26" => cos_16 <= x"AAEB" ;
        when x"A27" => cos_16 <= x"AB11" ;
        when x"A28" => cos_16 <= x"AB37" ;
        when x"A29" => cos_16 <= x"AB5C" ;
        when x"A2A" => cos_16 <= x"AB82" ;
        when x"A2B" => cos_16 <= x"ABA8" ;
        when x"A2C" => cos_16 <= x"ABCE" ;
        when x"A2D" => cos_16 <= x"ABF4" ;
        when x"A2E" => cos_16 <= x"AC19" ;
        when x"A2F" => cos_16 <= x"AC3F" ;
        when x"A30" => cos_16 <= x"AC65" ;
        when x"A31" => cos_16 <= x"AC8C" ;
        when x"A32" => cos_16 <= x"ACB2" ;
        when x"A33" => cos_16 <= x"ACD8" ;
        when x"A34" => cos_16 <= x"ACFE" ;
        when x"A35" => cos_16 <= x"AD24" ;
        when x"A36" => cos_16 <= x"AD4B" ;
        when x"A37" => cos_16 <= x"AD71" ;
        when x"A38" => cos_16 <= x"AD98" ;
        when x"A39" => cos_16 <= x"ADBE" ;
        when x"A3A" => cos_16 <= x"ADE5" ;
        when x"A3B" => cos_16 <= x"AE0B" ;
        when x"A3C" => cos_16 <= x"AE32" ;
        when x"A3D" => cos_16 <= x"AE58" ;
        when x"A3E" => cos_16 <= x"AE7F" ;
        when x"A3F" => cos_16 <= x"AEA6" ;
        when x"A40" => cos_16 <= x"AECD" ;
        when x"A41" => cos_16 <= x"AEF4" ;
        when x"A42" => cos_16 <= x"AF1B" ;
        when x"A43" => cos_16 <= x"AF42" ;
        when x"A44" => cos_16 <= x"AF69" ;
        when x"A45" => cos_16 <= x"AF90" ;
        when x"A46" => cos_16 <= x"AFB7" ;
        when x"A47" => cos_16 <= x"AFDE" ;
        when x"A48" => cos_16 <= x"B005" ;
        when x"A49" => cos_16 <= x"B02C" ;
        when x"A4A" => cos_16 <= x"B054" ;
        when x"A4B" => cos_16 <= x"B07B" ;
        when x"A4C" => cos_16 <= x"B0A3" ;
        when x"A4D" => cos_16 <= x"B0CA" ;
        when x"A4E" => cos_16 <= x"B0F2" ;
        when x"A4F" => cos_16 <= x"B119" ;
        when x"A50" => cos_16 <= x"B141" ;
        when x"A51" => cos_16 <= x"B168" ;
        when x"A52" => cos_16 <= x"B190" ;
        when x"A53" => cos_16 <= x"B1B8" ;
        when x"A54" => cos_16 <= x"B1E0" ;
        when x"A55" => cos_16 <= x"B207" ;
        when x"A56" => cos_16 <= x"B22F" ;
        when x"A57" => cos_16 <= x"B257" ;
        when x"A58" => cos_16 <= x"B27F" ;
        when x"A59" => cos_16 <= x"B2A7" ;
        when x"A5A" => cos_16 <= x"B2CF" ;
        when x"A5B" => cos_16 <= x"B2F7" ;
        when x"A5C" => cos_16 <= x"B320" ;
        when x"A5D" => cos_16 <= x"B348" ;
        when x"A5E" => cos_16 <= x"B370" ;
        when x"A5F" => cos_16 <= x"B398" ;
        when x"A60" => cos_16 <= x"B3C1" ;
        when x"A61" => cos_16 <= x"B3E9" ;
        when x"A62" => cos_16 <= x"B412" ;
        when x"A63" => cos_16 <= x"B43A" ;
        when x"A64" => cos_16 <= x"B463" ;
        when x"A65" => cos_16 <= x"B48B" ;
        when x"A66" => cos_16 <= x"B4B4" ;
        when x"A67" => cos_16 <= x"B4DC" ;
        when x"A68" => cos_16 <= x"B505" ;
        when x"A69" => cos_16 <= x"B52E" ;
        when x"A6A" => cos_16 <= x"B557" ;
        when x"A6B" => cos_16 <= x"B580" ;
        when x"A6C" => cos_16 <= x"B5A8" ;
        when x"A6D" => cos_16 <= x"B5D1" ;
        when x"A6E" => cos_16 <= x"B5FA" ;
        when x"A6F" => cos_16 <= x"B623" ;
        when x"A70" => cos_16 <= x"B64C" ;
        when x"A71" => cos_16 <= x"B676" ;
        when x"A72" => cos_16 <= x"B69F" ;
        when x"A73" => cos_16 <= x"B6C8" ;
        when x"A74" => cos_16 <= x"B6F1" ;
        when x"A75" => cos_16 <= x"B71B" ;
        when x"A76" => cos_16 <= x"B744" ;
        when x"A77" => cos_16 <= x"B76D" ;
        when x"A78" => cos_16 <= x"B797" ;
        when x"A79" => cos_16 <= x"B7C0" ;
        when x"A7A" => cos_16 <= x"B7EA" ;
        when x"A7B" => cos_16 <= x"B813" ;
        when x"A7C" => cos_16 <= x"B83D" ;
        when x"A7D" => cos_16 <= x"B866" ;
        when x"A7E" => cos_16 <= x"B890" ;
        when x"A7F" => cos_16 <= x"B8BA" ;
        when x"A80" => cos_16 <= x"B8E4" ;
        when x"A81" => cos_16 <= x"B90D" ;
        when x"A82" => cos_16 <= x"B937" ;
        when x"A83" => cos_16 <= x"B961" ;
        when x"A84" => cos_16 <= x"B98B" ;
        when x"A85" => cos_16 <= x"B9B5" ;
        when x"A86" => cos_16 <= x"B9DF" ;
        when x"A87" => cos_16 <= x"BA09" ;
        when x"A88" => cos_16 <= x"BA33" ;
        when x"A89" => cos_16 <= x"BA5D" ;
        when x"A8A" => cos_16 <= x"BA88" ;
        when x"A8B" => cos_16 <= x"BAB2" ;
        when x"A8C" => cos_16 <= x"BADC" ;
        when x"A8D" => cos_16 <= x"BB07" ;
        when x"A8E" => cos_16 <= x"BB31" ;
        when x"A8F" => cos_16 <= x"BB5B" ;
        when x"A90" => cos_16 <= x"BB86" ;
        when x"A91" => cos_16 <= x"BBB0" ;
        when x"A92" => cos_16 <= x"BBDB" ;
        when x"A93" => cos_16 <= x"BC05" ;
        when x"A94" => cos_16 <= x"BC30" ;
        when x"A95" => cos_16 <= x"BC5B" ;
        when x"A96" => cos_16 <= x"BC85" ;
        when x"A97" => cos_16 <= x"BCB0" ;
        when x"A98" => cos_16 <= x"BCDB" ;
        when x"A99" => cos_16 <= x"BD06" ;
        when x"A9A" => cos_16 <= x"BD30" ;
        when x"A9B" => cos_16 <= x"BD5B" ;
        when x"A9C" => cos_16 <= x"BD86" ;
        when x"A9D" => cos_16 <= x"BDB1" ;
        when x"A9E" => cos_16 <= x"BDDC" ;
        when x"A9F" => cos_16 <= x"BE07" ;
        when x"AA0" => cos_16 <= x"BE32" ;
        when x"AA1" => cos_16 <= x"BE5E" ;
        when x"AA2" => cos_16 <= x"BE89" ;
        when x"AA3" => cos_16 <= x"BEB4" ;
        when x"AA4" => cos_16 <= x"BEDF" ;
        when x"AA5" => cos_16 <= x"BF0A" ;
        when x"AA6" => cos_16 <= x"BF36" ;
        when x"AA7" => cos_16 <= x"BF61" ;
        when x"AA8" => cos_16 <= x"BF8D" ;
        when x"AA9" => cos_16 <= x"BFB8" ;
        when x"AAA" => cos_16 <= x"BFE3" ;
        when x"AAB" => cos_16 <= x"C00F" ;
        when x"AAC" => cos_16 <= x"C03B" ;
        when x"AAD" => cos_16 <= x"C066" ;
        when x"AAE" => cos_16 <= x"C092" ;
        when x"AAF" => cos_16 <= x"C0BD" ;
        when x"AB0" => cos_16 <= x"C0E9" ;
        when x"AB1" => cos_16 <= x"C115" ;
        when x"AB2" => cos_16 <= x"C141" ;
        when x"AB3" => cos_16 <= x"C16D" ;
        when x"AB4" => cos_16 <= x"C198" ;
        when x"AB5" => cos_16 <= x"C1C4" ;
        when x"AB6" => cos_16 <= x"C1F0" ;
        when x"AB7" => cos_16 <= x"C21C" ;
        when x"AB8" => cos_16 <= x"C248" ;
        when x"AB9" => cos_16 <= x"C274" ;
        when x"ABA" => cos_16 <= x"C2A0" ;
        when x"ABB" => cos_16 <= x"C2CD" ;
        when x"ABC" => cos_16 <= x"C2F9" ;
        when x"ABD" => cos_16 <= x"C325" ;
        when x"ABE" => cos_16 <= x"C351" ;
        when x"ABF" => cos_16 <= x"C37D" ;
        when x"AC0" => cos_16 <= x"C3AA" ;
        when x"AC1" => cos_16 <= x"C3D6" ;
        when x"AC2" => cos_16 <= x"C402" ;
        when x"AC3" => cos_16 <= x"C42F" ;
        when x"AC4" => cos_16 <= x"C45B" ;
        when x"AC5" => cos_16 <= x"C488" ;
        when x"AC6" => cos_16 <= x"C4B4" ;
        when x"AC7" => cos_16 <= x"C4E1" ;
        when x"AC8" => cos_16 <= x"C50E" ;
        when x"AC9" => cos_16 <= x"C53A" ;
        when x"ACA" => cos_16 <= x"C567" ;
        when x"ACB" => cos_16 <= x"C594" ;
        when x"ACC" => cos_16 <= x"C5C0" ;
        when x"ACD" => cos_16 <= x"C5ED" ;
        when x"ACE" => cos_16 <= x"C61A" ;
        when x"ACF" => cos_16 <= x"C647" ;
        when x"AD0" => cos_16 <= x"C674" ;
        when x"AD1" => cos_16 <= x"C6A0" ;
        when x"AD2" => cos_16 <= x"C6CD" ;
        when x"AD3" => cos_16 <= x"C6FA" ;
        when x"AD4" => cos_16 <= x"C727" ;
        when x"AD5" => cos_16 <= x"C755" ;
        when x"AD6" => cos_16 <= x"C782" ;
        when x"AD7" => cos_16 <= x"C7AF" ;
        when x"AD8" => cos_16 <= x"C7DC" ;
        when x"AD9" => cos_16 <= x"C809" ;
        when x"ADA" => cos_16 <= x"C836" ;
        when x"ADB" => cos_16 <= x"C864" ;
        when x"ADC" => cos_16 <= x"C891" ;
        when x"ADD" => cos_16 <= x"C8BE" ;
        when x"ADE" => cos_16 <= x"C8EB" ;
        when x"ADF" => cos_16 <= x"C919" ;
        when x"AE0" => cos_16 <= x"C946" ;
        when x"AE1" => cos_16 <= x"C974" ;
        when x"AE2" => cos_16 <= x"C9A1" ;
        when x"AE3" => cos_16 <= x"C9CF" ;
        when x"AE4" => cos_16 <= x"C9FC" ;
        when x"AE5" => cos_16 <= x"CA2A" ;
        when x"AE6" => cos_16 <= x"CA58" ;
        when x"AE7" => cos_16 <= x"CA85" ;
        when x"AE8" => cos_16 <= x"CAB3" ;
        when x"AE9" => cos_16 <= x"CAE1" ;
        when x"AEA" => cos_16 <= x"CB0E" ;
        when x"AEB" => cos_16 <= x"CB3C" ;
        when x"AEC" => cos_16 <= x"CB6A" ;
        when x"AED" => cos_16 <= x"CB98" ;
        when x"AEE" => cos_16 <= x"CBC6" ;
        when x"AEF" => cos_16 <= x"CBF4" ;
        when x"AF0" => cos_16 <= x"CC21" ;
        when x"AF1" => cos_16 <= x"CC4F" ;
        when x"AF2" => cos_16 <= x"CC7D" ;
        when x"AF3" => cos_16 <= x"CCAB" ;
        when x"AF4" => cos_16 <= x"CCDA" ;
        when x"AF5" => cos_16 <= x"CD08" ;
        when x"AF6" => cos_16 <= x"CD36" ;
        when x"AF7" => cos_16 <= x"CD64" ;
        when x"AF8" => cos_16 <= x"CD92" ;
        when x"AF9" => cos_16 <= x"CDC0" ;
        when x"AFA" => cos_16 <= x"CDEF" ;
        when x"AFB" => cos_16 <= x"CE1D" ;
        when x"AFC" => cos_16 <= x"CE4B" ;
        when x"AFD" => cos_16 <= x"CE79" ;
        when x"AFE" => cos_16 <= x"CEA8" ;
        when x"AFF" => cos_16 <= x"CED6" ;
        when x"B00" => cos_16 <= x"CF05" ;
        when x"B01" => cos_16 <= x"CF33" ;
        when x"B02" => cos_16 <= x"CF62" ;
        when x"B03" => cos_16 <= x"CF90" ;
        when x"B04" => cos_16 <= x"CFBF" ;
        when x"B05" => cos_16 <= x"CFED" ;
        when x"B06" => cos_16 <= x"D01C" ;
        when x"B07" => cos_16 <= x"D04A" ;
        when x"B08" => cos_16 <= x"D079" ;
        when x"B09" => cos_16 <= x"D0A8" ;
        when x"B0A" => cos_16 <= x"D0D6" ;
        when x"B0B" => cos_16 <= x"D105" ;
        when x"B0C" => cos_16 <= x"D134" ;
        when x"B0D" => cos_16 <= x"D163" ;
        when x"B0E" => cos_16 <= x"D192" ;
        when x"B0F" => cos_16 <= x"D1C0" ;
        when x"B10" => cos_16 <= x"D1EF" ;
        when x"B11" => cos_16 <= x"D21E" ;
        when x"B12" => cos_16 <= x"D24D" ;
        when x"B13" => cos_16 <= x"D27C" ;
        when x"B14" => cos_16 <= x"D2AB" ;
        when x"B15" => cos_16 <= x"D2DA" ;
        when x"B16" => cos_16 <= x"D309" ;
        when x"B17" => cos_16 <= x"D338" ;
        when x"B18" => cos_16 <= x"D367" ;
        when x"B19" => cos_16 <= x"D396" ;
        when x"B1A" => cos_16 <= x"D3C6" ;
        when x"B1B" => cos_16 <= x"D3F5" ;
        when x"B1C" => cos_16 <= x"D424" ;
        when x"B1D" => cos_16 <= x"D453" ;
        when x"B1E" => cos_16 <= x"D483" ;
        when x"B1F" => cos_16 <= x"D4B2" ;
        when x"B20" => cos_16 <= x"D4E1" ;
        when x"B21" => cos_16 <= x"D510" ;
        when x"B22" => cos_16 <= x"D540" ;
        when x"B23" => cos_16 <= x"D56F" ;
        when x"B24" => cos_16 <= x"D59F" ;
        when x"B25" => cos_16 <= x"D5CE" ;
        when x"B26" => cos_16 <= x"D5FE" ;
        when x"B27" => cos_16 <= x"D62D" ;
        when x"B28" => cos_16 <= x"D65D" ;
        when x"B29" => cos_16 <= x"D68C" ;
        when x"B2A" => cos_16 <= x"D6BC" ;
        when x"B2B" => cos_16 <= x"D6EB" ;
        when x"B2C" => cos_16 <= x"D71B" ;
        when x"B2D" => cos_16 <= x"D74B" ;
        when x"B2E" => cos_16 <= x"D77A" ;
        when x"B2F" => cos_16 <= x"D7AA" ;
        when x"B30" => cos_16 <= x"D7DA" ;
        when x"B31" => cos_16 <= x"D809" ;
        when x"B32" => cos_16 <= x"D839" ;
        when x"B33" => cos_16 <= x"D869" ;
        when x"B34" => cos_16 <= x"D899" ;
        when x"B35" => cos_16 <= x"D8C9" ;
        when x"B36" => cos_16 <= x"D8F8" ;
        when x"B37" => cos_16 <= x"D928" ;
        when x"B38" => cos_16 <= x"D958" ;
        when x"B39" => cos_16 <= x"D988" ;
        when x"B3A" => cos_16 <= x"D9B8" ;
        when x"B3B" => cos_16 <= x"D9E8" ;
        when x"B3C" => cos_16 <= x"DA18" ;
        when x"B3D" => cos_16 <= x"DA48" ;
        when x"B3E" => cos_16 <= x"DA78" ;
        when x"B3F" => cos_16 <= x"DAA8" ;
        when x"B40" => cos_16 <= x"DAD8" ;
        when x"B41" => cos_16 <= x"DB08" ;
        when x"B42" => cos_16 <= x"DB38" ;
        when x"B43" => cos_16 <= x"DB69" ;
        when x"B44" => cos_16 <= x"DB99" ;
        when x"B45" => cos_16 <= x"DBC9" ;
        when x"B46" => cos_16 <= x"DBF9" ;
        when x"B47" => cos_16 <= x"DC29" ;
        when x"B48" => cos_16 <= x"DC5A" ;
        when x"B49" => cos_16 <= x"DC8A" ;
        when x"B4A" => cos_16 <= x"DCBA" ;
        when x"B4B" => cos_16 <= x"DCEB" ;
        when x"B4C" => cos_16 <= x"DD1B" ;
        when x"B4D" => cos_16 <= x"DD4B" ;
        when x"B4E" => cos_16 <= x"DD7C" ;
        when x"B4F" => cos_16 <= x"DDAC" ;
        when x"B50" => cos_16 <= x"DDDD" ;
        when x"B51" => cos_16 <= x"DE0D" ;
        when x"B52" => cos_16 <= x"DE3E" ;
        when x"B53" => cos_16 <= x"DE6E" ;
        when x"B54" => cos_16 <= x"DE9F" ;
        when x"B55" => cos_16 <= x"DECF" ;
        when x"B56" => cos_16 <= x"DF00" ;
        when x"B57" => cos_16 <= x"DF30" ;
        when x"B58" => cos_16 <= x"DF61" ;
        when x"B59" => cos_16 <= x"DF91" ;
        when x"B5A" => cos_16 <= x"DFC2" ;
        when x"B5B" => cos_16 <= x"DFF3" ;
        when x"B5C" => cos_16 <= x"E023" ;
        when x"B5D" => cos_16 <= x"E054" ;
        when x"B5E" => cos_16 <= x"E085" ;
        when x"B5F" => cos_16 <= x"E0B6" ;
        when x"B60" => cos_16 <= x"E0E6" ;
        when x"B61" => cos_16 <= x"E117" ;
        when x"B62" => cos_16 <= x"E148" ;
        when x"B63" => cos_16 <= x"E179" ;
        when x"B64" => cos_16 <= x"E1A9" ;
        when x"B65" => cos_16 <= x"E1DA" ;
        when x"B66" => cos_16 <= x"E20B" ;
        when x"B67" => cos_16 <= x"E23C" ;
        when x"B68" => cos_16 <= x"E26D" ;
        when x"B69" => cos_16 <= x"E29E" ;
        when x"B6A" => cos_16 <= x"E2CF" ;
        when x"B6B" => cos_16 <= x"E300" ;
        when x"B6C" => cos_16 <= x"E331" ;
        when x"B6D" => cos_16 <= x"E362" ;
        when x"B6E" => cos_16 <= x"E393" ;
        when x"B6F" => cos_16 <= x"E3C4" ;
        when x"B70" => cos_16 <= x"E3F5" ;
        when x"B71" => cos_16 <= x"E426" ;
        when x"B72" => cos_16 <= x"E457" ;
        when x"B73" => cos_16 <= x"E488" ;
        when x"B74" => cos_16 <= x"E4B9" ;
        when x"B75" => cos_16 <= x"E4EA" ;
        when x"B76" => cos_16 <= x"E51B" ;
        when x"B77" => cos_16 <= x"E54C" ;
        when x"B78" => cos_16 <= x"E57E" ;
        when x"B79" => cos_16 <= x"E5AF" ;
        when x"B7A" => cos_16 <= x"E5E0" ;
        when x"B7B" => cos_16 <= x"E611" ;
        when x"B7C" => cos_16 <= x"E642" ;
        when x"B7D" => cos_16 <= x"E674" ;
        when x"B7E" => cos_16 <= x"E6A5" ;
        when x"B7F" => cos_16 <= x"E6D6" ;
        when x"B80" => cos_16 <= x"E707" ;
        when x"B81" => cos_16 <= x"E739" ;
        when x"B82" => cos_16 <= x"E76A" ;
        when x"B83" => cos_16 <= x"E79B" ;
        when x"B84" => cos_16 <= x"E7CD" ;
        when x"B85" => cos_16 <= x"E7FE" ;
        when x"B86" => cos_16 <= x"E830" ;
        when x"B87" => cos_16 <= x"E861" ;
        when x"B88" => cos_16 <= x"E892" ;
        when x"B89" => cos_16 <= x"E8C4" ;
        when x"B8A" => cos_16 <= x"E8F5" ;
        when x"B8B" => cos_16 <= x"E927" ;
        when x"B8C" => cos_16 <= x"E958" ;
        when x"B8D" => cos_16 <= x"E98A" ;
        when x"B8E" => cos_16 <= x"E9BB" ;
        when x"B8F" => cos_16 <= x"E9ED" ;
        when x"B90" => cos_16 <= x"EA1E" ;
        when x"B91" => cos_16 <= x"EA50" ;
        when x"B92" => cos_16 <= x"EA81" ;
        when x"B93" => cos_16 <= x"EAB3" ;
        when x"B94" => cos_16 <= x"EAE4" ;
        when x"B95" => cos_16 <= x"EB16" ;
        when x"B96" => cos_16 <= x"EB47" ;
        when x"B97" => cos_16 <= x"EB79" ;
        when x"B98" => cos_16 <= x"EBAB" ;
        when x"B99" => cos_16 <= x"EBDC" ;
        when x"B9A" => cos_16 <= x"EC0E" ;
        when x"B9B" => cos_16 <= x"EC40" ;
        when x"B9C" => cos_16 <= x"EC71" ;
        when x"B9D" => cos_16 <= x"ECA3" ;
        when x"B9E" => cos_16 <= x"ECD5" ;
        when x"B9F" => cos_16 <= x"ED06" ;
        when x"BA0" => cos_16 <= x"ED38" ;
        when x"BA1" => cos_16 <= x"ED6A" ;
        when x"BA2" => cos_16 <= x"ED9C" ;
        when x"BA3" => cos_16 <= x"EDCD" ;
        when x"BA4" => cos_16 <= x"EDFF" ;
        when x"BA5" => cos_16 <= x"EE31" ;
        when x"BA6" => cos_16 <= x"EE63" ;
        when x"BA7" => cos_16 <= x"EE94" ;
        when x"BA8" => cos_16 <= x"EEC6" ;
        when x"BA9" => cos_16 <= x"EEF8" ;
        when x"BAA" => cos_16 <= x"EF2A" ;
        when x"BAB" => cos_16 <= x"EF5C" ;
        when x"BAC" => cos_16 <= x"EF8E" ;
        when x"BAD" => cos_16 <= x"EFBF" ;
        when x"BAE" => cos_16 <= x"EFF1" ;
        when x"BAF" => cos_16 <= x"F023" ;
        when x"BB0" => cos_16 <= x"F055" ;
        when x"BB1" => cos_16 <= x"F087" ;
        when x"BB2" => cos_16 <= x"F0B9" ;
        when x"BB3" => cos_16 <= x"F0EB" ;
        when x"BB4" => cos_16 <= x"F11D" ;
        when x"BB5" => cos_16 <= x"F14F" ;
        when x"BB6" => cos_16 <= x"F180" ;
        when x"BB7" => cos_16 <= x"F1B2" ;
        when x"BB8" => cos_16 <= x"F1E4" ;
        when x"BB9" => cos_16 <= x"F216" ;
        when x"BBA" => cos_16 <= x"F248" ;
        when x"BBB" => cos_16 <= x"F27A" ;
        when x"BBC" => cos_16 <= x"F2AC" ;
        when x"BBD" => cos_16 <= x"F2DE" ;
        when x"BBE" => cos_16 <= x"F310" ;
        when x"BBF" => cos_16 <= x"F342" ;
        when x"BC0" => cos_16 <= x"F374" ;
        when x"BC1" => cos_16 <= x"F3A6" ;
        when x"BC2" => cos_16 <= x"F3D8" ;
        when x"BC3" => cos_16 <= x"F40A" ;
        when x"BC4" => cos_16 <= x"F43C" ;
        when x"BC5" => cos_16 <= x"F46E" ;
        when x"BC6" => cos_16 <= x"F4A1" ;
        when x"BC7" => cos_16 <= x"F4D3" ;
        when x"BC8" => cos_16 <= x"F505" ;
        when x"BC9" => cos_16 <= x"F537" ;
        when x"BCA" => cos_16 <= x"F569" ;
        when x"BCB" => cos_16 <= x"F59B" ;
        when x"BCC" => cos_16 <= x"F5CD" ;
        when x"BCD" => cos_16 <= x"F5FF" ;
        when x"BCE" => cos_16 <= x"F631" ;
        when x"BCF" => cos_16 <= x"F663" ;
        when x"BD0" => cos_16 <= x"F696" ;
        when x"BD1" => cos_16 <= x"F6C8" ;
        when x"BD2" => cos_16 <= x"F6FA" ;
        when x"BD3" => cos_16 <= x"F72C" ;
        when x"BD4" => cos_16 <= x"F75E" ;
        when x"BD5" => cos_16 <= x"F790" ;
        when x"BD6" => cos_16 <= x"F7C2" ;
        when x"BD7" => cos_16 <= x"F7F5" ;
        when x"BD8" => cos_16 <= x"F827" ;
        when x"BD9" => cos_16 <= x"F859" ;
        when x"BDA" => cos_16 <= x"F88B" ;
        when x"BDB" => cos_16 <= x"F8BD" ;
        when x"BDC" => cos_16 <= x"F8EF" ;
        when x"BDD" => cos_16 <= x"F922" ;
        when x"BDE" => cos_16 <= x"F954" ;
        when x"BDF" => cos_16 <= x"F986" ;
        when x"BE0" => cos_16 <= x"F9B8" ;
        when x"BE1" => cos_16 <= x"F9EA" ;
        when x"BE2" => cos_16 <= x"FA1D" ;
        when x"BE3" => cos_16 <= x"FA4F" ;
        when x"BE4" => cos_16 <= x"FA81" ;
        when x"BE5" => cos_16 <= x"FAB3" ;
        when x"BE6" => cos_16 <= x"FAE5" ;
        when x"BE7" => cos_16 <= x"FB18" ;
        when x"BE8" => cos_16 <= x"FB4A" ;
        when x"BE9" => cos_16 <= x"FB7C" ;
        when x"BEA" => cos_16 <= x"FBAE" ;
        when x"BEB" => cos_16 <= x"FBE1" ;
        when x"BEC" => cos_16 <= x"FC13" ;
        when x"BED" => cos_16 <= x"FC45" ;
        when x"BEE" => cos_16 <= x"FC77" ;
        when x"BEF" => cos_16 <= x"FCAA" ;
        when x"BF0" => cos_16 <= x"FCDC" ;
        when x"BF1" => cos_16 <= x"FD0E" ;
        when x"BF2" => cos_16 <= x"FD40" ;
        when x"BF3" => cos_16 <= x"FD73" ;
        when x"BF4" => cos_16 <= x"FDA5" ;
        when x"BF5" => cos_16 <= x"FDD7" ;
        when x"BF6" => cos_16 <= x"FE09" ;
        when x"BF7" => cos_16 <= x"FE3C" ;
        when x"BF8" => cos_16 <= x"FE6E" ;
        when x"BF9" => cos_16 <= x"FEA0" ;
        when x"BFA" => cos_16 <= x"FED2" ;
        when x"BFB" => cos_16 <= x"FF05" ;
        when x"BFC" => cos_16 <= x"FF37" ;
        when x"BFD" => cos_16 <= x"FF69" ;
        when x"BFE" => cos_16 <= x"FF9B" ;
        when x"BFF" => cos_16 <= x"FFCE" ;
        when x"C00" => cos_16 <= x"0000" ;
        when x"C01" => cos_16 <= x"0032" ;
        when x"C02" => cos_16 <= x"0065" ;
        when x"C03" => cos_16 <= x"0097" ;
        when x"C04" => cos_16 <= x"00C9" ;
        when x"C05" => cos_16 <= x"00FB" ;
        when x"C06" => cos_16 <= x"012E" ;
        when x"C07" => cos_16 <= x"0160" ;
        when x"C08" => cos_16 <= x"0192" ;
        when x"C09" => cos_16 <= x"01C4" ;
        when x"C0A" => cos_16 <= x"01F7" ;
        when x"C0B" => cos_16 <= x"0229" ;
        when x"C0C" => cos_16 <= x"025B" ;
        when x"C0D" => cos_16 <= x"028D" ;
        when x"C0E" => cos_16 <= x"02C0" ;
        when x"C0F" => cos_16 <= x"02F2" ;
        when x"C10" => cos_16 <= x"0324" ;
        when x"C11" => cos_16 <= x"0356" ;
        when x"C12" => cos_16 <= x"0389" ;
        when x"C13" => cos_16 <= x"03BB" ;
        when x"C14" => cos_16 <= x"03ED" ;
        when x"C15" => cos_16 <= x"041F" ;
        when x"C16" => cos_16 <= x"0452" ;
        when x"C17" => cos_16 <= x"0484" ;
        when x"C18" => cos_16 <= x"04B6" ;
        when x"C19" => cos_16 <= x"04E8" ;
        when x"C1A" => cos_16 <= x"051B" ;
        when x"C1B" => cos_16 <= x"054D" ;
        when x"C1C" => cos_16 <= x"057F" ;
        when x"C1D" => cos_16 <= x"05B1" ;
        when x"C1E" => cos_16 <= x"05E3" ;
        when x"C1F" => cos_16 <= x"0616" ;
        when x"C20" => cos_16 <= x"0648" ;
        when x"C21" => cos_16 <= x"067A" ;
        when x"C22" => cos_16 <= x"06AC" ;
        when x"C23" => cos_16 <= x"06DE" ;
        when x"C24" => cos_16 <= x"0711" ;
        when x"C25" => cos_16 <= x"0743" ;
        when x"C26" => cos_16 <= x"0775" ;
        when x"C27" => cos_16 <= x"07A7" ;
        when x"C28" => cos_16 <= x"07D9" ;
        when x"C29" => cos_16 <= x"080B" ;
        when x"C2A" => cos_16 <= x"083E" ;
        when x"C2B" => cos_16 <= x"0870" ;
        when x"C2C" => cos_16 <= x"08A2" ;
        when x"C2D" => cos_16 <= x"08D4" ;
        when x"C2E" => cos_16 <= x"0906" ;
        when x"C2F" => cos_16 <= x"0938" ;
        when x"C30" => cos_16 <= x"096A" ;
        when x"C31" => cos_16 <= x"099D" ;
        when x"C32" => cos_16 <= x"09CF" ;
        when x"C33" => cos_16 <= x"0A01" ;
        when x"C34" => cos_16 <= x"0A33" ;
        when x"C35" => cos_16 <= x"0A65" ;
        when x"C36" => cos_16 <= x"0A97" ;
        when x"C37" => cos_16 <= x"0AC9" ;
        when x"C38" => cos_16 <= x"0AFB" ;
        when x"C39" => cos_16 <= x"0B2D" ;
        when x"C3A" => cos_16 <= x"0B5F" ;
        when x"C3B" => cos_16 <= x"0B92" ;
        when x"C3C" => cos_16 <= x"0BC4" ;
        when x"C3D" => cos_16 <= x"0BF6" ;
        when x"C3E" => cos_16 <= x"0C28" ;
        when x"C3F" => cos_16 <= x"0C5A" ;
        when x"C40" => cos_16 <= x"0C8C" ;
        when x"C41" => cos_16 <= x"0CBE" ;
        when x"C42" => cos_16 <= x"0CF0" ;
        when x"C43" => cos_16 <= x"0D22" ;
        when x"C44" => cos_16 <= x"0D54" ;
        when x"C45" => cos_16 <= x"0D86" ;
        when x"C46" => cos_16 <= x"0DB8" ;
        when x"C47" => cos_16 <= x"0DEA" ;
        when x"C48" => cos_16 <= x"0E1C" ;
        when x"C49" => cos_16 <= x"0E4E" ;
        when x"C4A" => cos_16 <= x"0E80" ;
        when x"C4B" => cos_16 <= x"0EB1" ;
        when x"C4C" => cos_16 <= x"0EE3" ;
        when x"C4D" => cos_16 <= x"0F15" ;
        when x"C4E" => cos_16 <= x"0F47" ;
        when x"C4F" => cos_16 <= x"0F79" ;
        when x"C50" => cos_16 <= x"0FAB" ;
        when x"C51" => cos_16 <= x"0FDD" ;
        when x"C52" => cos_16 <= x"100F" ;
        when x"C53" => cos_16 <= x"1041" ;
        when x"C54" => cos_16 <= x"1072" ;
        when x"C55" => cos_16 <= x"10A4" ;
        when x"C56" => cos_16 <= x"10D6" ;
        when x"C57" => cos_16 <= x"1108" ;
        when x"C58" => cos_16 <= x"113A" ;
        when x"C59" => cos_16 <= x"116C" ;
        when x"C5A" => cos_16 <= x"119D" ;
        when x"C5B" => cos_16 <= x"11CF" ;
        when x"C5C" => cos_16 <= x"1201" ;
        when x"C5D" => cos_16 <= x"1233" ;
        when x"C5E" => cos_16 <= x"1264" ;
        when x"C5F" => cos_16 <= x"1296" ;
        when x"C60" => cos_16 <= x"12C8" ;
        when x"C61" => cos_16 <= x"12FA" ;
        when x"C62" => cos_16 <= x"132B" ;
        when x"C63" => cos_16 <= x"135D" ;
        when x"C64" => cos_16 <= x"138F" ;
        when x"C65" => cos_16 <= x"13C0" ;
        when x"C66" => cos_16 <= x"13F2" ;
        when x"C67" => cos_16 <= x"1424" ;
        when x"C68" => cos_16 <= x"1455" ;
        when x"C69" => cos_16 <= x"1487" ;
        when x"C6A" => cos_16 <= x"14B9" ;
        when x"C6B" => cos_16 <= x"14EA" ;
        when x"C6C" => cos_16 <= x"151C" ;
        when x"C6D" => cos_16 <= x"154D" ;
        when x"C6E" => cos_16 <= x"157F" ;
        when x"C6F" => cos_16 <= x"15B0" ;
        when x"C70" => cos_16 <= x"15E2" ;
        when x"C71" => cos_16 <= x"1613" ;
        when x"C72" => cos_16 <= x"1645" ;
        when x"C73" => cos_16 <= x"1676" ;
        when x"C74" => cos_16 <= x"16A8" ;
        when x"C75" => cos_16 <= x"16D9" ;
        when x"C76" => cos_16 <= x"170B" ;
        when x"C77" => cos_16 <= x"173C" ;
        when x"C78" => cos_16 <= x"176E" ;
        when x"C79" => cos_16 <= x"179F" ;
        when x"C7A" => cos_16 <= x"17D0" ;
        when x"C7B" => cos_16 <= x"1802" ;
        when x"C7C" => cos_16 <= x"1833" ;
        when x"C7D" => cos_16 <= x"1865" ;
        when x"C7E" => cos_16 <= x"1896" ;
        when x"C7F" => cos_16 <= x"18C7" ;
        when x"C80" => cos_16 <= x"18F9" ;
        when x"C81" => cos_16 <= x"192A" ;
        when x"C82" => cos_16 <= x"195B" ;
        when x"C83" => cos_16 <= x"198C" ;
        when x"C84" => cos_16 <= x"19BE" ;
        when x"C85" => cos_16 <= x"19EF" ;
        when x"C86" => cos_16 <= x"1A20" ;
        when x"C87" => cos_16 <= x"1A51" ;
        when x"C88" => cos_16 <= x"1A82" ;
        when x"C89" => cos_16 <= x"1AB4" ;
        when x"C8A" => cos_16 <= x"1AE5" ;
        when x"C8B" => cos_16 <= x"1B16" ;
        when x"C8C" => cos_16 <= x"1B47" ;
        when x"C8D" => cos_16 <= x"1B78" ;
        when x"C8E" => cos_16 <= x"1BA9" ;
        when x"C8F" => cos_16 <= x"1BDA" ;
        when x"C90" => cos_16 <= x"1C0B" ;
        when x"C91" => cos_16 <= x"1C3C" ;
        when x"C92" => cos_16 <= x"1C6D" ;
        when x"C93" => cos_16 <= x"1C9E" ;
        when x"C94" => cos_16 <= x"1CCF" ;
        when x"C95" => cos_16 <= x"1D00" ;
        when x"C96" => cos_16 <= x"1D31" ;
        when x"C97" => cos_16 <= x"1D62" ;
        when x"C98" => cos_16 <= x"1D93" ;
        when x"C99" => cos_16 <= x"1DC4" ;
        when x"C9A" => cos_16 <= x"1DF5" ;
        when x"C9B" => cos_16 <= x"1E26" ;
        when x"C9C" => cos_16 <= x"1E57" ;
        when x"C9D" => cos_16 <= x"1E87" ;
        when x"C9E" => cos_16 <= x"1EB8" ;
        when x"C9F" => cos_16 <= x"1EE9" ;
        when x"CA0" => cos_16 <= x"1F1A" ;
        when x"CA1" => cos_16 <= x"1F4A" ;
        when x"CA2" => cos_16 <= x"1F7B" ;
        when x"CA3" => cos_16 <= x"1FAC" ;
        when x"CA4" => cos_16 <= x"1FDD" ;
        when x"CA5" => cos_16 <= x"200D" ;
        when x"CA6" => cos_16 <= x"203E" ;
        when x"CA7" => cos_16 <= x"206F" ;
        when x"CA8" => cos_16 <= x"209F" ;
        when x"CA9" => cos_16 <= x"20D0" ;
        when x"CAA" => cos_16 <= x"2100" ;
        when x"CAB" => cos_16 <= x"2131" ;
        when x"CAC" => cos_16 <= x"2161" ;
        when x"CAD" => cos_16 <= x"2192" ;
        when x"CAE" => cos_16 <= x"21C2" ;
        when x"CAF" => cos_16 <= x"21F3" ;
        when x"CB0" => cos_16 <= x"2223" ;
        when x"CB1" => cos_16 <= x"2254" ;
        when x"CB2" => cos_16 <= x"2284" ;
        when x"CB3" => cos_16 <= x"22B5" ;
        when x"CB4" => cos_16 <= x"22E5" ;
        when x"CB5" => cos_16 <= x"2315" ;
        when x"CB6" => cos_16 <= x"2346" ;
        when x"CB7" => cos_16 <= x"2376" ;
        when x"CB8" => cos_16 <= x"23A6" ;
        when x"CB9" => cos_16 <= x"23D7" ;
        when x"CBA" => cos_16 <= x"2407" ;
        when x"CBB" => cos_16 <= x"2437" ;
        when x"CBC" => cos_16 <= x"2467" ;
        when x"CBD" => cos_16 <= x"2497" ;
        when x"CBE" => cos_16 <= x"24C8" ;
        when x"CBF" => cos_16 <= x"24F8" ;
        when x"CC0" => cos_16 <= x"2528" ;
        when x"CC1" => cos_16 <= x"2558" ;
        when x"CC2" => cos_16 <= x"2588" ;
        when x"CC3" => cos_16 <= x"25B8" ;
        when x"CC4" => cos_16 <= x"25E8" ;
        when x"CC5" => cos_16 <= x"2618" ;
        when x"CC6" => cos_16 <= x"2648" ;
        when x"CC7" => cos_16 <= x"2678" ;
        when x"CC8" => cos_16 <= x"26A8" ;
        when x"CC9" => cos_16 <= x"26D8" ;
        when x"CCA" => cos_16 <= x"2708" ;
        when x"CCB" => cos_16 <= x"2737" ;
        when x"CCC" => cos_16 <= x"2767" ;
        when x"CCD" => cos_16 <= x"2797" ;
        when x"CCE" => cos_16 <= x"27C7" ;
        when x"CCF" => cos_16 <= x"27F7" ;
        when x"CD0" => cos_16 <= x"2826" ;
        when x"CD1" => cos_16 <= x"2856" ;
        when x"CD2" => cos_16 <= x"2886" ;
        when x"CD3" => cos_16 <= x"28B5" ;
        when x"CD4" => cos_16 <= x"28E5" ;
        when x"CD5" => cos_16 <= x"2915" ;
        when x"CD6" => cos_16 <= x"2944" ;
        when x"CD7" => cos_16 <= x"2974" ;
        when x"CD8" => cos_16 <= x"29A3" ;
        when x"CD9" => cos_16 <= x"29D3" ;
        when x"CDA" => cos_16 <= x"2A02" ;
        when x"CDB" => cos_16 <= x"2A32" ;
        when x"CDC" => cos_16 <= x"2A61" ;
        when x"CDD" => cos_16 <= x"2A91" ;
        when x"CDE" => cos_16 <= x"2AC0" ;
        when x"CDF" => cos_16 <= x"2AF0" ;
        when x"CE0" => cos_16 <= x"2B1F" ;
        when x"CE1" => cos_16 <= x"2B4E" ;
        when x"CE2" => cos_16 <= x"2B7D" ;
        when x"CE3" => cos_16 <= x"2BAD" ;
        when x"CE4" => cos_16 <= x"2BDC" ;
        when x"CE5" => cos_16 <= x"2C0B" ;
        when x"CE6" => cos_16 <= x"2C3A" ;
        when x"CE7" => cos_16 <= x"2C6A" ;
        when x"CE8" => cos_16 <= x"2C99" ;
        when x"CE9" => cos_16 <= x"2CC8" ;
        when x"CEA" => cos_16 <= x"2CF7" ;
        when x"CEB" => cos_16 <= x"2D26" ;
        when x"CEC" => cos_16 <= x"2D55" ;
        when x"CED" => cos_16 <= x"2D84" ;
        when x"CEE" => cos_16 <= x"2DB3" ;
        when x"CEF" => cos_16 <= x"2DE2" ;
        when x"CF0" => cos_16 <= x"2E11" ;
        when x"CF1" => cos_16 <= x"2E40" ;
        when x"CF2" => cos_16 <= x"2E6E" ;
        when x"CF3" => cos_16 <= x"2E9D" ;
        when x"CF4" => cos_16 <= x"2ECC" ;
        when x"CF5" => cos_16 <= x"2EFB" ;
        when x"CF6" => cos_16 <= x"2F2A" ;
        when x"CF7" => cos_16 <= x"2F58" ;
        when x"CF8" => cos_16 <= x"2F87" ;
        when x"CF9" => cos_16 <= x"2FB6" ;
        when x"CFA" => cos_16 <= x"2FE4" ;
        when x"CFB" => cos_16 <= x"3013" ;
        when x"CFC" => cos_16 <= x"3041" ;
        when x"CFD" => cos_16 <= x"3070" ;
        when x"CFE" => cos_16 <= x"309E" ;
        when x"CFF" => cos_16 <= x"30CD" ;
        when x"D00" => cos_16 <= x"30FB" ;
        when x"D01" => cos_16 <= x"312A" ;
        when x"D02" => cos_16 <= x"3158" ;
        when x"D03" => cos_16 <= x"3187" ;
        when x"D04" => cos_16 <= x"31B5" ;
        when x"D05" => cos_16 <= x"31E3" ;
        when x"D06" => cos_16 <= x"3211" ;
        when x"D07" => cos_16 <= x"3240" ;
        when x"D08" => cos_16 <= x"326E" ;
        when x"D09" => cos_16 <= x"329C" ;
        when x"D0A" => cos_16 <= x"32CA" ;
        when x"D0B" => cos_16 <= x"32F8" ;
        when x"D0C" => cos_16 <= x"3326" ;
        when x"D0D" => cos_16 <= x"3355" ;
        when x"D0E" => cos_16 <= x"3383" ;
        when x"D0F" => cos_16 <= x"33B1" ;
        when x"D10" => cos_16 <= x"33DF" ;
        when x"D11" => cos_16 <= x"340C" ;
        when x"D12" => cos_16 <= x"343A" ;
        when x"D13" => cos_16 <= x"3468" ;
        when x"D14" => cos_16 <= x"3496" ;
        when x"D15" => cos_16 <= x"34C4" ;
        when x"D16" => cos_16 <= x"34F2" ;
        when x"D17" => cos_16 <= x"351F" ;
        when x"D18" => cos_16 <= x"354D" ;
        when x"D19" => cos_16 <= x"357B" ;
        when x"D1A" => cos_16 <= x"35A8" ;
        when x"D1B" => cos_16 <= x"35D6" ;
        when x"D1C" => cos_16 <= x"3604" ;
        when x"D1D" => cos_16 <= x"3631" ;
        when x"D1E" => cos_16 <= x"365F" ;
        when x"D1F" => cos_16 <= x"368C" ;
        when x"D20" => cos_16 <= x"36BA" ;
        when x"D21" => cos_16 <= x"36E7" ;
        when x"D22" => cos_16 <= x"3715" ;
        when x"D23" => cos_16 <= x"3742" ;
        when x"D24" => cos_16 <= x"376F" ;
        when x"D25" => cos_16 <= x"379C" ;
        when x"D26" => cos_16 <= x"37CA" ;
        when x"D27" => cos_16 <= x"37F7" ;
        when x"D28" => cos_16 <= x"3824" ;
        when x"D29" => cos_16 <= x"3851" ;
        when x"D2A" => cos_16 <= x"387E" ;
        when x"D2B" => cos_16 <= x"38AB" ;
        when x"D2C" => cos_16 <= x"38D9" ;
        when x"D2D" => cos_16 <= x"3906" ;
        when x"D2E" => cos_16 <= x"3933" ;
        when x"D2F" => cos_16 <= x"3960" ;
        when x"D30" => cos_16 <= x"398C" ;
        when x"D31" => cos_16 <= x"39B9" ;
        when x"D32" => cos_16 <= x"39E6" ;
        when x"D33" => cos_16 <= x"3A13" ;
        when x"D34" => cos_16 <= x"3A40" ;
        when x"D35" => cos_16 <= x"3A6C" ;
        when x"D36" => cos_16 <= x"3A99" ;
        when x"D37" => cos_16 <= x"3AC6" ;
        when x"D38" => cos_16 <= x"3AF2" ;
        when x"D39" => cos_16 <= x"3B1F" ;
        when x"D3A" => cos_16 <= x"3B4C" ;
        when x"D3B" => cos_16 <= x"3B78" ;
        when x"D3C" => cos_16 <= x"3BA5" ;
        when x"D3D" => cos_16 <= x"3BD1" ;
        when x"D3E" => cos_16 <= x"3BFE" ;
        when x"D3F" => cos_16 <= x"3C2A" ;
        when x"D40" => cos_16 <= x"3C56" ;
        when x"D41" => cos_16 <= x"3C83" ;
        when x"D42" => cos_16 <= x"3CAF" ;
        when x"D43" => cos_16 <= x"3CDB" ;
        when x"D44" => cos_16 <= x"3D07" ;
        when x"D45" => cos_16 <= x"3D33" ;
        when x"D46" => cos_16 <= x"3D60" ;
        when x"D47" => cos_16 <= x"3D8C" ;
        when x"D48" => cos_16 <= x"3DB8" ;
        when x"D49" => cos_16 <= x"3DE4" ;
        when x"D4A" => cos_16 <= x"3E10" ;
        when x"D4B" => cos_16 <= x"3E3C" ;
        when x"D4C" => cos_16 <= x"3E68" ;
        when x"D4D" => cos_16 <= x"3E93" ;
        when x"D4E" => cos_16 <= x"3EBF" ;
        when x"D4F" => cos_16 <= x"3EEB" ;
        when x"D50" => cos_16 <= x"3F17" ;
        when x"D51" => cos_16 <= x"3F43" ;
        when x"D52" => cos_16 <= x"3F6E" ;
        when x"D53" => cos_16 <= x"3F9A" ;
        when x"D54" => cos_16 <= x"3FC5" ;
        when x"D55" => cos_16 <= x"3FF1" ;
        when x"D56" => cos_16 <= x"401D" ;
        when x"D57" => cos_16 <= x"4048" ;
        when x"D58" => cos_16 <= x"4073" ;
        when x"D59" => cos_16 <= x"409F" ;
        when x"D5A" => cos_16 <= x"40CA" ;
        when x"D5B" => cos_16 <= x"40F6" ;
        when x"D5C" => cos_16 <= x"4121" ;
        when x"D5D" => cos_16 <= x"414C" ;
        when x"D5E" => cos_16 <= x"4177" ;
        when x"D5F" => cos_16 <= x"41A2" ;
        when x"D60" => cos_16 <= x"41CE" ;
        when x"D61" => cos_16 <= x"41F9" ;
        when x"D62" => cos_16 <= x"4224" ;
        when x"D63" => cos_16 <= x"424F" ;
        when x"D64" => cos_16 <= x"427A" ;
        when x"D65" => cos_16 <= x"42A5" ;
        when x"D66" => cos_16 <= x"42D0" ;
        when x"D67" => cos_16 <= x"42FA" ;
        when x"D68" => cos_16 <= x"4325" ;
        when x"D69" => cos_16 <= x"4350" ;
        when x"D6A" => cos_16 <= x"437B" ;
        when x"D6B" => cos_16 <= x"43A5" ;
        when x"D6C" => cos_16 <= x"43D0" ;
        when x"D6D" => cos_16 <= x"43FB" ;
        when x"D6E" => cos_16 <= x"4425" ;
        when x"D6F" => cos_16 <= x"4450" ;
        when x"D70" => cos_16 <= x"447A" ;
        when x"D71" => cos_16 <= x"44A5" ;
        when x"D72" => cos_16 <= x"44CF" ;
        when x"D73" => cos_16 <= x"44F9" ;
        when x"D74" => cos_16 <= x"4524" ;
        when x"D75" => cos_16 <= x"454E" ;
        when x"D76" => cos_16 <= x"4578" ;
        when x"D77" => cos_16 <= x"45A3" ;
        when x"D78" => cos_16 <= x"45CD" ;
        when x"D79" => cos_16 <= x"45F7" ;
        when x"D7A" => cos_16 <= x"4621" ;
        when x"D7B" => cos_16 <= x"464B" ;
        when x"D7C" => cos_16 <= x"4675" ;
        when x"D7D" => cos_16 <= x"469F" ;
        when x"D7E" => cos_16 <= x"46C9" ;
        when x"D7F" => cos_16 <= x"46F3" ;
        when x"D80" => cos_16 <= x"471C" ;
        when x"D81" => cos_16 <= x"4746" ;
        when x"D82" => cos_16 <= x"4770" ;
        when x"D83" => cos_16 <= x"479A" ;
        when x"D84" => cos_16 <= x"47C3" ;
        when x"D85" => cos_16 <= x"47ED" ;
        when x"D86" => cos_16 <= x"4816" ;
        when x"D87" => cos_16 <= x"4840" ;
        when x"D88" => cos_16 <= x"4869" ;
        when x"D89" => cos_16 <= x"4893" ;
        when x"D8A" => cos_16 <= x"48BC" ;
        when x"D8B" => cos_16 <= x"48E5" ;
        when x"D8C" => cos_16 <= x"490F" ;
        when x"D8D" => cos_16 <= x"4938" ;
        when x"D8E" => cos_16 <= x"4961" ;
        when x"D8F" => cos_16 <= x"498A" ;
        when x"D90" => cos_16 <= x"49B4" ;
        when x"D91" => cos_16 <= x"49DD" ;
        when x"D92" => cos_16 <= x"4A06" ;
        when x"D93" => cos_16 <= x"4A2F" ;
        when x"D94" => cos_16 <= x"4A58" ;
        when x"D95" => cos_16 <= x"4A80" ;
        when x"D96" => cos_16 <= x"4AA9" ;
        when x"D97" => cos_16 <= x"4AD2" ;
        when x"D98" => cos_16 <= x"4AFB" ;
        when x"D99" => cos_16 <= x"4B24" ;
        when x"D9A" => cos_16 <= x"4B4C" ;
        when x"D9B" => cos_16 <= x"4B75" ;
        when x"D9C" => cos_16 <= x"4B9D" ;
        when x"D9D" => cos_16 <= x"4BC6" ;
        when x"D9E" => cos_16 <= x"4BEE" ;
        when x"D9F" => cos_16 <= x"4C17" ;
        when x"DA0" => cos_16 <= x"4C3F" ;
        when x"DA1" => cos_16 <= x"4C68" ;
        when x"DA2" => cos_16 <= x"4C90" ;
        when x"DA3" => cos_16 <= x"4CB8" ;
        when x"DA4" => cos_16 <= x"4CE0" ;
        when x"DA5" => cos_16 <= x"4D09" ;
        when x"DA6" => cos_16 <= x"4D31" ;
        when x"DA7" => cos_16 <= x"4D59" ;
        when x"DA8" => cos_16 <= x"4D81" ;
        when x"DA9" => cos_16 <= x"4DA9" ;
        when x"DAA" => cos_16 <= x"4DD1" ;
        when x"DAB" => cos_16 <= x"4DF9" ;
        when x"DAC" => cos_16 <= x"4E20" ;
        when x"DAD" => cos_16 <= x"4E48" ;
        when x"DAE" => cos_16 <= x"4E70" ;
        when x"DAF" => cos_16 <= x"4E98" ;
        when x"DB0" => cos_16 <= x"4EBF" ;
        when x"DB1" => cos_16 <= x"4EE7" ;
        when x"DB2" => cos_16 <= x"4F0E" ;
        when x"DB3" => cos_16 <= x"4F36" ;
        when x"DB4" => cos_16 <= x"4F5D" ;
        when x"DB5" => cos_16 <= x"4F85" ;
        when x"DB6" => cos_16 <= x"4FAC" ;
        when x"DB7" => cos_16 <= x"4FD4" ;
        when x"DB8" => cos_16 <= x"4FFB" ;
        when x"DB9" => cos_16 <= x"5022" ;
        when x"DBA" => cos_16 <= x"5049" ;
        when x"DBB" => cos_16 <= x"5070" ;
        when x"DBC" => cos_16 <= x"5097" ;
        when x"DBD" => cos_16 <= x"50BE" ;
        when x"DBE" => cos_16 <= x"50E5" ;
        when x"DBF" => cos_16 <= x"510C" ;
        when x"DC0" => cos_16 <= x"5133" ;
        when x"DC1" => cos_16 <= x"515A" ;
        when x"DC2" => cos_16 <= x"5181" ;
        when x"DC3" => cos_16 <= x"51A8" ;
        when x"DC4" => cos_16 <= x"51CE" ;
        when x"DC5" => cos_16 <= x"51F5" ;
        when x"DC6" => cos_16 <= x"521B" ;
        when x"DC7" => cos_16 <= x"5242" ;
        when x"DC8" => cos_16 <= x"5268" ;
        when x"DC9" => cos_16 <= x"528F" ;
        when x"DCA" => cos_16 <= x"52B5" ;
        when x"DCB" => cos_16 <= x"52DC" ;
        when x"DCC" => cos_16 <= x"5302" ;
        when x"DCD" => cos_16 <= x"5328" ;
        when x"DCE" => cos_16 <= x"534E" ;
        when x"DCF" => cos_16 <= x"5374" ;
        when x"DD0" => cos_16 <= x"539B" ;
        when x"DD1" => cos_16 <= x"53C1" ;
        when x"DD2" => cos_16 <= x"53E7" ;
        when x"DD3" => cos_16 <= x"540C" ;
        when x"DD4" => cos_16 <= x"5432" ;
        when x"DD5" => cos_16 <= x"5458" ;
        when x"DD6" => cos_16 <= x"547E" ;
        when x"DD7" => cos_16 <= x"54A4" ;
        when x"DD8" => cos_16 <= x"54C9" ;
        when x"DD9" => cos_16 <= x"54EF" ;
        when x"DDA" => cos_16 <= x"5515" ;
        when x"DDB" => cos_16 <= x"553A" ;
        when x"DDC" => cos_16 <= x"5560" ;
        when x"DDD" => cos_16 <= x"5585" ;
        when x"DDE" => cos_16 <= x"55AA" ;
        when x"DDF" => cos_16 <= x"55D0" ;
        when x"DE0" => cos_16 <= x"55F5" ;
        when x"DE1" => cos_16 <= x"561A" ;
        when x"DE2" => cos_16 <= x"563F" ;
        when x"DE3" => cos_16 <= x"5664" ;
        when x"DE4" => cos_16 <= x"568A" ;
        when x"DE5" => cos_16 <= x"56AF" ;
        when x"DE6" => cos_16 <= x"56D3" ;
        when x"DE7" => cos_16 <= x"56F8" ;
        when x"DE8" => cos_16 <= x"571D" ;
        when x"DE9" => cos_16 <= x"5742" ;
        when x"DEA" => cos_16 <= x"5767" ;
        when x"DEB" => cos_16 <= x"578B" ;
        when x"DEC" => cos_16 <= x"57B0" ;
        when x"DED" => cos_16 <= x"57D5" ;
        when x"DEE" => cos_16 <= x"57F9" ;
        when x"DEF" => cos_16 <= x"581E" ;
        when x"DF0" => cos_16 <= x"5842" ;
        when x"DF1" => cos_16 <= x"5867" ;
        when x"DF2" => cos_16 <= x"588B" ;
        when x"DF3" => cos_16 <= x"58AF" ;
        when x"DF4" => cos_16 <= x"58D3" ;
        when x"DF5" => cos_16 <= x"58F8" ;
        when x"DF6" => cos_16 <= x"591C" ;
        when x"DF7" => cos_16 <= x"5940" ;
        when x"DF8" => cos_16 <= x"5964" ;
        when x"DF9" => cos_16 <= x"5988" ;
        when x"DFA" => cos_16 <= x"59AC" ;
        when x"DFB" => cos_16 <= x"59CF" ;
        when x"DFC" => cos_16 <= x"59F3" ;
        when x"DFD" => cos_16 <= x"5A17" ;
        when x"DFE" => cos_16 <= x"5A3B" ;
        when x"DFF" => cos_16 <= x"5A5E" ;
        when x"E00" => cos_16 <= x"5A82" ;
        when x"E01" => cos_16 <= x"5AA5" ;
        when x"E02" => cos_16 <= x"5AC9" ;
        when x"E03" => cos_16 <= x"5AEC" ;
        when x"E04" => cos_16 <= x"5B0F" ;
        when x"E05" => cos_16 <= x"5B33" ;
        when x"E06" => cos_16 <= x"5B56" ;
        when x"E07" => cos_16 <= x"5B79" ;
        when x"E08" => cos_16 <= x"5B9C" ;
        when x"E09" => cos_16 <= x"5BBF" ;
        when x"E0A" => cos_16 <= x"5BE2" ;
        when x"E0B" => cos_16 <= x"5C05" ;
        when x"E0C" => cos_16 <= x"5C28" ;
        when x"E0D" => cos_16 <= x"5C4B" ;
        when x"E0E" => cos_16 <= x"5C6E" ;
        when x"E0F" => cos_16 <= x"5C91" ;
        when x"E10" => cos_16 <= x"5CB3" ;
        when x"E11" => cos_16 <= x"5CD6" ;
        when x"E12" => cos_16 <= x"5CF9" ;
        when x"E13" => cos_16 <= x"5D1B" ;
        when x"E14" => cos_16 <= x"5D3E" ;
        when x"E15" => cos_16 <= x"5D60" ;
        when x"E16" => cos_16 <= x"5D82" ;
        when x"E17" => cos_16 <= x"5DA5" ;
        when x"E18" => cos_16 <= x"5DC7" ;
        when x"E19" => cos_16 <= x"5DE9" ;
        when x"E1A" => cos_16 <= x"5E0B" ;
        when x"E1B" => cos_16 <= x"5E2D" ;
        when x"E1C" => cos_16 <= x"5E4F" ;
        when x"E1D" => cos_16 <= x"5E71" ;
        when x"E1E" => cos_16 <= x"5E93" ;
        when x"E1F" => cos_16 <= x"5EB5" ;
        when x"E20" => cos_16 <= x"5ED7" ;
        when x"E21" => cos_16 <= x"5EF8" ;
        when x"E22" => cos_16 <= x"5F1A" ;
        when x"E23" => cos_16 <= x"5F3C" ;
        when x"E24" => cos_16 <= x"5F5D" ;
        when x"E25" => cos_16 <= x"5F7F" ;
        when x"E26" => cos_16 <= x"5FA0" ;
        when x"E27" => cos_16 <= x"5FC2" ;
        when x"E28" => cos_16 <= x"5FE3" ;
        when x"E29" => cos_16 <= x"6004" ;
        when x"E2A" => cos_16 <= x"6025" ;
        when x"E2B" => cos_16 <= x"6047" ;
        when x"E2C" => cos_16 <= x"6068" ;
        when x"E2D" => cos_16 <= x"6089" ;
        when x"E2E" => cos_16 <= x"60AA" ;
        when x"E2F" => cos_16 <= x"60CB" ;
        when x"E30" => cos_16 <= x"60EB" ;
        when x"E31" => cos_16 <= x"610C" ;
        when x"E32" => cos_16 <= x"612D" ;
        when x"E33" => cos_16 <= x"614E" ;
        when x"E34" => cos_16 <= x"616E" ;
        when x"E35" => cos_16 <= x"618F" ;
        when x"E36" => cos_16 <= x"61AF" ;
        when x"E37" => cos_16 <= x"61D0" ;
        when x"E38" => cos_16 <= x"61F0" ;
        when x"E39" => cos_16 <= x"6211" ;
        when x"E3A" => cos_16 <= x"6231" ;
        when x"E3B" => cos_16 <= x"6251" ;
        when x"E3C" => cos_16 <= x"6271" ;
        when x"E3D" => cos_16 <= x"6291" ;
        when x"E3E" => cos_16 <= x"62B1" ;
        when x"E3F" => cos_16 <= x"62D1" ;
        when x"E40" => cos_16 <= x"62F1" ;
        when x"E41" => cos_16 <= x"6311" ;
        when x"E42" => cos_16 <= x"6331" ;
        when x"E43" => cos_16 <= x"6351" ;
        when x"E44" => cos_16 <= x"6370" ;
        when x"E45" => cos_16 <= x"6390" ;
        when x"E46" => cos_16 <= x"63AF" ;
        when x"E47" => cos_16 <= x"63CF" ;
        when x"E48" => cos_16 <= x"63EE" ;
        when x"E49" => cos_16 <= x"640E" ;
        when x"E4A" => cos_16 <= x"642D" ;
        when x"E4B" => cos_16 <= x"644C" ;
        when x"E4C" => cos_16 <= x"646C" ;
        when x"E4D" => cos_16 <= x"648B" ;
        when x"E4E" => cos_16 <= x"64AA" ;
        when x"E4F" => cos_16 <= x"64C9" ;
        when x"E50" => cos_16 <= x"64E8" ;
        when x"E51" => cos_16 <= x"6507" ;
        when x"E52" => cos_16 <= x"6525" ;
        when x"E53" => cos_16 <= x"6544" ;
        when x"E54" => cos_16 <= x"6563" ;
        when x"E55" => cos_16 <= x"6582" ;
        when x"E56" => cos_16 <= x"65A0" ;
        when x"E57" => cos_16 <= x"65BF" ;
        when x"E58" => cos_16 <= x"65DD" ;
        when x"E59" => cos_16 <= x"65FC" ;
        when x"E5A" => cos_16 <= x"661A" ;
        when x"E5B" => cos_16 <= x"6638" ;
        when x"E5C" => cos_16 <= x"6656" ;
        when x"E5D" => cos_16 <= x"6675" ;
        when x"E5E" => cos_16 <= x"6693" ;
        when x"E5F" => cos_16 <= x"66B1" ;
        when x"E60" => cos_16 <= x"66CF" ;
        when x"E61" => cos_16 <= x"66ED" ;
        when x"E62" => cos_16 <= x"670A" ;
        when x"E63" => cos_16 <= x"6728" ;
        when x"E64" => cos_16 <= x"6746" ;
        when x"E65" => cos_16 <= x"6764" ;
        when x"E66" => cos_16 <= x"6781" ;
        when x"E67" => cos_16 <= x"679F" ;
        when x"E68" => cos_16 <= x"67BC" ;
        when x"E69" => cos_16 <= x"67DA" ;
        when x"E6A" => cos_16 <= x"67F7" ;
        when x"E6B" => cos_16 <= x"6814" ;
        when x"E6C" => cos_16 <= x"6832" ;
        when x"E6D" => cos_16 <= x"684F" ;
        when x"E6E" => cos_16 <= x"686C" ;
        when x"E6F" => cos_16 <= x"6889" ;
        when x"E70" => cos_16 <= x"68A6" ;
        when x"E71" => cos_16 <= x"68C3" ;
        when x"E72" => cos_16 <= x"68E0" ;
        when x"E73" => cos_16 <= x"68FC" ;
        when x"E74" => cos_16 <= x"6919" ;
        when x"E75" => cos_16 <= x"6936" ;
        when x"E76" => cos_16 <= x"6952" ;
        when x"E77" => cos_16 <= x"696F" ;
        when x"E78" => cos_16 <= x"698B" ;
        when x"E79" => cos_16 <= x"69A8" ;
        when x"E7A" => cos_16 <= x"69C4" ;
        when x"E7B" => cos_16 <= x"69E0" ;
        when x"E7C" => cos_16 <= x"69FD" ;
        when x"E7D" => cos_16 <= x"6A19" ;
        when x"E7E" => cos_16 <= x"6A35" ;
        when x"E7F" => cos_16 <= x"6A51" ;
        when x"E80" => cos_16 <= x"6A6D" ;
        when x"E81" => cos_16 <= x"6A89" ;
        when x"E82" => cos_16 <= x"6AA4" ;
        when x"E83" => cos_16 <= x"6AC0" ;
        when x"E84" => cos_16 <= x"6ADC" ;
        when x"E85" => cos_16 <= x"6AF8" ;
        when x"E86" => cos_16 <= x"6B13" ;
        when x"E87" => cos_16 <= x"6B2F" ;
        when x"E88" => cos_16 <= x"6B4A" ;
        when x"E89" => cos_16 <= x"6B65" ;
        when x"E8A" => cos_16 <= x"6B81" ;
        when x"E8B" => cos_16 <= x"6B9C" ;
        when x"E8C" => cos_16 <= x"6BB7" ;
        when x"E8D" => cos_16 <= x"6BD2" ;
        when x"E8E" => cos_16 <= x"6BED" ;
        when x"E8F" => cos_16 <= x"6C08" ;
        when x"E90" => cos_16 <= x"6C23" ;
        when x"E91" => cos_16 <= x"6C3E" ;
        when x"E92" => cos_16 <= x"6C59" ;
        when x"E93" => cos_16 <= x"6C74" ;
        when x"E94" => cos_16 <= x"6C8E" ;
        when x"E95" => cos_16 <= x"6CA9" ;
        when x"E96" => cos_16 <= x"6CC3" ;
        when x"E97" => cos_16 <= x"6CDE" ;
        when x"E98" => cos_16 <= x"6CF8" ;
        when x"E99" => cos_16 <= x"6D13" ;
        when x"E9A" => cos_16 <= x"6D2D" ;
        when x"E9B" => cos_16 <= x"6D47" ;
        when x"E9C" => cos_16 <= x"6D61" ;
        when x"E9D" => cos_16 <= x"6D7B" ;
        when x"E9E" => cos_16 <= x"6D95" ;
        when x"E9F" => cos_16 <= x"6DAF" ;
        when x"EA0" => cos_16 <= x"6DC9" ;
        when x"EA1" => cos_16 <= x"6DE3" ;
        when x"EA2" => cos_16 <= x"6DFD" ;
        when x"EA3" => cos_16 <= x"6E16" ;
        when x"EA4" => cos_16 <= x"6E30" ;
        when x"EA5" => cos_16 <= x"6E4A" ;
        when x"EA6" => cos_16 <= x"6E63" ;
        when x"EA7" => cos_16 <= x"6E7C" ;
        when x"EA8" => cos_16 <= x"6E96" ;
        when x"EA9" => cos_16 <= x"6EAF" ;
        when x"EAA" => cos_16 <= x"6EC8" ;
        when x"EAB" => cos_16 <= x"6EE1" ;
        when x"EAC" => cos_16 <= x"6EFB" ;
        when x"EAD" => cos_16 <= x"6F14" ;
        when x"EAE" => cos_16 <= x"6F2C" ;
        when x"EAF" => cos_16 <= x"6F45" ;
        when x"EB0" => cos_16 <= x"6F5E" ;
        when x"EB1" => cos_16 <= x"6F77" ;
        when x"EB2" => cos_16 <= x"6F90" ;
        when x"EB3" => cos_16 <= x"6FA8" ;
        when x"EB4" => cos_16 <= x"6FC1" ;
        when x"EB5" => cos_16 <= x"6FD9" ;
        when x"EB6" => cos_16 <= x"6FF2" ;
        when x"EB7" => cos_16 <= x"700A" ;
        when x"EB8" => cos_16 <= x"7022" ;
        when x"EB9" => cos_16 <= x"703A" ;
        when x"EBA" => cos_16 <= x"7053" ;
        when x"EBB" => cos_16 <= x"706B" ;
        when x"EBC" => cos_16 <= x"7083" ;
        when x"EBD" => cos_16 <= x"709B" ;
        when x"EBE" => cos_16 <= x"70B2" ;
        when x"EBF" => cos_16 <= x"70CA" ;
        when x"EC0" => cos_16 <= x"70E2" ;
        when x"EC1" => cos_16 <= x"70FA" ;
        when x"EC2" => cos_16 <= x"7111" ;
        when x"EC3" => cos_16 <= x"7129" ;
        when x"EC4" => cos_16 <= x"7140" ;
        when x"EC5" => cos_16 <= x"7158" ;
        when x"EC6" => cos_16 <= x"716F" ;
        when x"EC7" => cos_16 <= x"7186" ;
        when x"EC8" => cos_16 <= x"719D" ;
        when x"EC9" => cos_16 <= x"71B4" ;
        when x"ECA" => cos_16 <= x"71CB" ;
        when x"ECB" => cos_16 <= x"71E2" ;
        when x"ECC" => cos_16 <= x"71F9" ;
        when x"ECD" => cos_16 <= x"7210" ;
        when x"ECE" => cos_16 <= x"7227" ;
        when x"ECF" => cos_16 <= x"723E" ;
        when x"ED0" => cos_16 <= x"7254" ;
        when x"ED1" => cos_16 <= x"726B" ;
        when x"ED2" => cos_16 <= x"7281" ;
        when x"ED3" => cos_16 <= x"7298" ;
        when x"ED4" => cos_16 <= x"72AE" ;
        when x"ED5" => cos_16 <= x"72C4" ;
        when x"ED6" => cos_16 <= x"72DB" ;
        when x"ED7" => cos_16 <= x"72F1" ;
        when x"ED8" => cos_16 <= x"7307" ;
        when x"ED9" => cos_16 <= x"731D" ;
        when x"EDA" => cos_16 <= x"7333" ;
        when x"EDB" => cos_16 <= x"7349" ;
        when x"EDC" => cos_16 <= x"735E" ;
        when x"EDD" => cos_16 <= x"7374" ;
        when x"EDE" => cos_16 <= x"738A" ;
        when x"EDF" => cos_16 <= x"739F" ;
        when x"EE0" => cos_16 <= x"73B5" ;
        when x"EE1" => cos_16 <= x"73CA" ;
        when x"EE2" => cos_16 <= x"73E0" ;
        when x"EE3" => cos_16 <= x"73F5" ;
        when x"EE4" => cos_16 <= x"740A" ;
        when x"EE5" => cos_16 <= x"7420" ;
        when x"EE6" => cos_16 <= x"7435" ;
        when x"EE7" => cos_16 <= x"744A" ;
        when x"EE8" => cos_16 <= x"745F" ;
        when x"EE9" => cos_16 <= x"7474" ;
        when x"EEA" => cos_16 <= x"7488" ;
        when x"EEB" => cos_16 <= x"749D" ;
        when x"EEC" => cos_16 <= x"74B2" ;
        when x"EED" => cos_16 <= x"74C6" ;
        when x"EEE" => cos_16 <= x"74DB" ;
        when x"EEF" => cos_16 <= x"74F0" ;
        when x"EF0" => cos_16 <= x"7504" ;
        when x"EF1" => cos_16 <= x"7518" ;
        when x"EF2" => cos_16 <= x"752D" ;
        when x"EF3" => cos_16 <= x"7541" ;
        when x"EF4" => cos_16 <= x"7555" ;
        when x"EF5" => cos_16 <= x"7569" ;
        when x"EF6" => cos_16 <= x"757D" ;
        when x"EF7" => cos_16 <= x"7591" ;
        when x"EF8" => cos_16 <= x"75A5" ;
        when x"EF9" => cos_16 <= x"75B8" ;
        when x"EFA" => cos_16 <= x"75CC" ;
        when x"EFB" => cos_16 <= x"75E0" ;
        when x"EFC" => cos_16 <= x"75F3" ;
        when x"EFD" => cos_16 <= x"7607" ;
        when x"EFE" => cos_16 <= x"761A" ;
        when x"EFF" => cos_16 <= x"762D" ;
        when x"F00" => cos_16 <= x"7641" ;
        when x"F01" => cos_16 <= x"7654" ;
        when x"F02" => cos_16 <= x"7667" ;
        when x"F03" => cos_16 <= x"767A" ;
        when x"F04" => cos_16 <= x"768D" ;
        when x"F05" => cos_16 <= x"76A0" ;
        when x"F06" => cos_16 <= x"76B3" ;
        when x"F07" => cos_16 <= x"76C6" ;
        when x"F08" => cos_16 <= x"76D8" ;
        when x"F09" => cos_16 <= x"76EB" ;
        when x"F0A" => cos_16 <= x"76FE" ;
        when x"F0B" => cos_16 <= x"7710" ;
        when x"F0C" => cos_16 <= x"7722" ;
        when x"F0D" => cos_16 <= x"7735" ;
        when x"F0E" => cos_16 <= x"7747" ;
        when x"F0F" => cos_16 <= x"7759" ;
        when x"F10" => cos_16 <= x"776B" ;
        when x"F11" => cos_16 <= x"777D" ;
        when x"F12" => cos_16 <= x"778F" ;
        when x"F13" => cos_16 <= x"77A1" ;
        when x"F14" => cos_16 <= x"77B3" ;
        when x"F15" => cos_16 <= x"77C5" ;
        when x"F16" => cos_16 <= x"77D7" ;
        when x"F17" => cos_16 <= x"77E8" ;
        when x"F18" => cos_16 <= x"77FA" ;
        when x"F19" => cos_16 <= x"780B" ;
        when x"F1A" => cos_16 <= x"781D" ;
        when x"F1B" => cos_16 <= x"782E" ;
        when x"F1C" => cos_16 <= x"783F" ;
        when x"F1D" => cos_16 <= x"7850" ;
        when x"F1E" => cos_16 <= x"7862" ;
        when x"F1F" => cos_16 <= x"7873" ;
        when x"F20" => cos_16 <= x"7884" ;
        when x"F21" => cos_16 <= x"7894" ;
        when x"F22" => cos_16 <= x"78A5" ;
        when x"F23" => cos_16 <= x"78B6" ;
        when x"F24" => cos_16 <= x"78C7" ;
        when x"F25" => cos_16 <= x"78D7" ;
        when x"F26" => cos_16 <= x"78E8" ;
        when x"F27" => cos_16 <= x"78F8" ;
        when x"F28" => cos_16 <= x"7909" ;
        when x"F29" => cos_16 <= x"7919" ;
        when x"F2A" => cos_16 <= x"7929" ;
        when x"F2B" => cos_16 <= x"7939" ;
        when x"F2C" => cos_16 <= x"794A" ;
        when x"F2D" => cos_16 <= x"795A" ;
        when x"F2E" => cos_16 <= x"796A" ;
        when x"F2F" => cos_16 <= x"7979" ;
        when x"F30" => cos_16 <= x"7989" ;
        when x"F31" => cos_16 <= x"7999" ;
        when x"F32" => cos_16 <= x"79A9" ;
        when x"F33" => cos_16 <= x"79B8" ;
        when x"F34" => cos_16 <= x"79C8" ;
        when x"F35" => cos_16 <= x"79D7" ;
        when x"F36" => cos_16 <= x"79E6" ;
        when x"F37" => cos_16 <= x"79F6" ;
        when x"F38" => cos_16 <= x"7A05" ;
        when x"F39" => cos_16 <= x"7A14" ;
        when x"F3A" => cos_16 <= x"7A23" ;
        when x"F3B" => cos_16 <= x"7A32" ;
        when x"F3C" => cos_16 <= x"7A41" ;
        when x"F3D" => cos_16 <= x"7A50" ;
        when x"F3E" => cos_16 <= x"7A5F" ;
        when x"F3F" => cos_16 <= x"7A6D" ;
        when x"F40" => cos_16 <= x"7A7C" ;
        when x"F41" => cos_16 <= x"7A8B" ;
        when x"F42" => cos_16 <= x"7A99" ;
        when x"F43" => cos_16 <= x"7AA8" ;
        when x"F44" => cos_16 <= x"7AB6" ;
        when x"F45" => cos_16 <= x"7AC4" ;
        when x"F46" => cos_16 <= x"7AD2" ;
        when x"F47" => cos_16 <= x"7AE0" ;
        when x"F48" => cos_16 <= x"7AEE" ;
        when x"F49" => cos_16 <= x"7AFC" ;
        when x"F4A" => cos_16 <= x"7B0A" ;
        when x"F4B" => cos_16 <= x"7B18" ;
        when x"F4C" => cos_16 <= x"7B26" ;
        when x"F4D" => cos_16 <= x"7B33" ;
        when x"F4E" => cos_16 <= x"7B41" ;
        when x"F4F" => cos_16 <= x"7B4F" ;
        when x"F50" => cos_16 <= x"7B5C" ;
        when x"F51" => cos_16 <= x"7B69" ;
        when x"F52" => cos_16 <= x"7B77" ;
        when x"F53" => cos_16 <= x"7B84" ;
        when x"F54" => cos_16 <= x"7B91" ;
        when x"F55" => cos_16 <= x"7B9E" ;
        when x"F56" => cos_16 <= x"7BAB" ;
        when x"F57" => cos_16 <= x"7BB8" ;
        when x"F58" => cos_16 <= x"7BC5" ;
        when x"F59" => cos_16 <= x"7BD2" ;
        when x"F5A" => cos_16 <= x"7BDE" ;
        when x"F5B" => cos_16 <= x"7BEB" ;
        when x"F5C" => cos_16 <= x"7BF8" ;
        when x"F5D" => cos_16 <= x"7C04" ;
        when x"F5E" => cos_16 <= x"7C10" ;
        when x"F5F" => cos_16 <= x"7C1D" ;
        when x"F60" => cos_16 <= x"7C29" ;
        when x"F61" => cos_16 <= x"7C35" ;
        when x"F62" => cos_16 <= x"7C41" ;
        when x"F63" => cos_16 <= x"7C4D" ;
        when x"F64" => cos_16 <= x"7C59" ;
        when x"F65" => cos_16 <= x"7C65" ;
        when x"F66" => cos_16 <= x"7C71" ;
        when x"F67" => cos_16 <= x"7C7D" ;
        when x"F68" => cos_16 <= x"7C88" ;
        when x"F69" => cos_16 <= x"7C94" ;
        when x"F6A" => cos_16 <= x"7C9F" ;
        when x"F6B" => cos_16 <= x"7CAB" ;
        when x"F6C" => cos_16 <= x"7CB6" ;
        when x"F6D" => cos_16 <= x"7CC1" ;
        when x"F6E" => cos_16 <= x"7CCD" ;
        when x"F6F" => cos_16 <= x"7CD8" ;
        when x"F70" => cos_16 <= x"7CE3" ;
        when x"F71" => cos_16 <= x"7CEE" ;
        when x"F72" => cos_16 <= x"7CF9" ;
        when x"F73" => cos_16 <= x"7D04" ;
        when x"F74" => cos_16 <= x"7D0E" ;
        when x"F75" => cos_16 <= x"7D19" ;
        when x"F76" => cos_16 <= x"7D24" ;
        when x"F77" => cos_16 <= x"7D2E" ;
        when x"F78" => cos_16 <= x"7D39" ;
        when x"F79" => cos_16 <= x"7D43" ;
        when x"F7A" => cos_16 <= x"7D4D" ;
        when x"F7B" => cos_16 <= x"7D57" ;
        when x"F7C" => cos_16 <= x"7D62" ;
        when x"F7D" => cos_16 <= x"7D6C" ;
        when x"F7E" => cos_16 <= x"7D76" ;
        when x"F7F" => cos_16 <= x"7D80" ;
        when x"F80" => cos_16 <= x"7D89" ;
        when x"F81" => cos_16 <= x"7D93" ;
        when x"F82" => cos_16 <= x"7D9D" ;
        when x"F83" => cos_16 <= x"7DA6" ;
        when x"F84" => cos_16 <= x"7DB0" ;
        when x"F85" => cos_16 <= x"7DB9" ;
        when x"F86" => cos_16 <= x"7DC3" ;
        when x"F87" => cos_16 <= x"7DCC" ;
        when x"F88" => cos_16 <= x"7DD5" ;
        when x"F89" => cos_16 <= x"7DDF" ;
        when x"F8A" => cos_16 <= x"7DE8" ;
        when x"F8B" => cos_16 <= x"7DF1" ;
        when x"F8C" => cos_16 <= x"7DFA" ;
        when x"F8D" => cos_16 <= x"7E02" ;
        when x"F8E" => cos_16 <= x"7E0B" ;
        when x"F8F" => cos_16 <= x"7E14" ;
        when x"F90" => cos_16 <= x"7E1D" ;
        when x"F91" => cos_16 <= x"7E25" ;
        when x"F92" => cos_16 <= x"7E2E" ;
        when x"F93" => cos_16 <= x"7E36" ;
        when x"F94" => cos_16 <= x"7E3E" ;
        when x"F95" => cos_16 <= x"7E47" ;
        when x"F96" => cos_16 <= x"7E4F" ;
        when x"F97" => cos_16 <= x"7E57" ;
        when x"F98" => cos_16 <= x"7E5F" ;
        when x"F99" => cos_16 <= x"7E67" ;
        when x"F9A" => cos_16 <= x"7E6F" ;
        when x"F9B" => cos_16 <= x"7E77" ;
        when x"F9C" => cos_16 <= x"7E7E" ;
        when x"F9D" => cos_16 <= x"7E86" ;
        when x"F9E" => cos_16 <= x"7E8D" ;
        when x"F9F" => cos_16 <= x"7E95" ;
        when x"FA0" => cos_16 <= x"7E9C" ;
        when x"FA1" => cos_16 <= x"7EA4" ;
        when x"FA2" => cos_16 <= x"7EAB" ;
        when x"FA3" => cos_16 <= x"7EB2" ;
        when x"FA4" => cos_16 <= x"7EB9" ;
        when x"FA5" => cos_16 <= x"7EC0" ;
        when x"FA6" => cos_16 <= x"7EC7" ;
        when x"FA7" => cos_16 <= x"7ECE" ;
        when x"FA8" => cos_16 <= x"7ED5" ;
        when x"FA9" => cos_16 <= x"7EDC" ;
        when x"FAA" => cos_16 <= x"7EE2" ;
        when x"FAB" => cos_16 <= x"7EE9" ;
        when x"FAC" => cos_16 <= x"7EEF" ;
        when x"FAD" => cos_16 <= x"7EF6" ;
        when x"FAE" => cos_16 <= x"7EFC" ;
        when x"FAF" => cos_16 <= x"7F02" ;
        when x"FB0" => cos_16 <= x"7F09" ;
        when x"FB1" => cos_16 <= x"7F0F" ;
        when x"FB2" => cos_16 <= x"7F15" ;
        when x"FB3" => cos_16 <= x"7F1B" ;
        when x"FB4" => cos_16 <= x"7F21" ;
        when x"FB5" => cos_16 <= x"7F26" ;
        when x"FB6" => cos_16 <= x"7F2C" ;
        when x"FB7" => cos_16 <= x"7F32" ;
        when x"FB8" => cos_16 <= x"7F37" ;
        when x"FB9" => cos_16 <= x"7F3D" ;
        when x"FBA" => cos_16 <= x"7F42" ;
        when x"FBB" => cos_16 <= x"7F48" ;
        when x"FBC" => cos_16 <= x"7F4D" ;
        when x"FBD" => cos_16 <= x"7F52" ;
        when x"FBE" => cos_16 <= x"7F57" ;
        when x"FBF" => cos_16 <= x"7F5C" ;
        when x"FC0" => cos_16 <= x"7F61" ;
        when x"FC1" => cos_16 <= x"7F66" ;
        when x"FC2" => cos_16 <= x"7F6B" ;
        when x"FC3" => cos_16 <= x"7F70" ;
        when x"FC4" => cos_16 <= x"7F74" ;
        when x"FC5" => cos_16 <= x"7F79" ;
        when x"FC6" => cos_16 <= x"7F7D" ;
        when x"FC7" => cos_16 <= x"7F82" ;
        when x"FC8" => cos_16 <= x"7F86" ;
        when x"FC9" => cos_16 <= x"7F8A" ;
        when x"FCA" => cos_16 <= x"7F8F" ;
        when x"FCB" => cos_16 <= x"7F93" ;
        when x"FCC" => cos_16 <= x"7F97" ;
        when x"FCD" => cos_16 <= x"7F9B" ;
        when x"FCE" => cos_16 <= x"7F9F" ;
        when x"FCF" => cos_16 <= x"7FA2" ;
        when x"FD0" => cos_16 <= x"7FA6" ;
        when x"FD1" => cos_16 <= x"7FAA" ;
        when x"FD2" => cos_16 <= x"7FAD" ;
        when x"FD3" => cos_16 <= x"7FB1" ;
        when x"FD4" => cos_16 <= x"7FB4" ;
        when x"FD5" => cos_16 <= x"7FB8" ;
        when x"FD6" => cos_16 <= x"7FBB" ;
        when x"FD7" => cos_16 <= x"7FBE" ;
        when x"FD8" => cos_16 <= x"7FC1" ;
        when x"FD9" => cos_16 <= x"7FC4" ;
        when x"FDA" => cos_16 <= x"7FC7" ;
        when x"FDB" => cos_16 <= x"7FCA" ;
        when x"FDC" => cos_16 <= x"7FCD" ;
        when x"FDD" => cos_16 <= x"7FD0" ;
        when x"FDE" => cos_16 <= x"7FD2" ;
        when x"FDF" => cos_16 <= x"7FD5" ;
        when x"FE0" => cos_16 <= x"7FD8" ;
        when x"FE1" => cos_16 <= x"7FDA" ;
        when x"FE2" => cos_16 <= x"7FDC" ;
        when x"FE3" => cos_16 <= x"7FDF" ;
        when x"FE4" => cos_16 <= x"7FE1" ;
        when x"FE5" => cos_16 <= x"7FE3" ;
        when x"FE6" => cos_16 <= x"7FE5" ;
        when x"FE7" => cos_16 <= x"7FE7" ;
        when x"FE8" => cos_16 <= x"7FE9" ;
        when x"FE9" => cos_16 <= x"7FEB" ;
        when x"FEA" => cos_16 <= x"7FEC" ;
        when x"FEB" => cos_16 <= x"7FEE" ;
        when x"FEC" => cos_16 <= x"7FF0" ;
        when x"FED" => cos_16 <= x"7FF1" ;
        when x"FEE" => cos_16 <= x"7FF3" ;
        when x"FEF" => cos_16 <= x"7FF4" ;
        when x"FF0" => cos_16 <= x"7FF5" ;
        when x"FF1" => cos_16 <= x"7FF6" ;
        when x"FF2" => cos_16 <= x"7FF7" ;
        when x"FF3" => cos_16 <= x"7FF8" ;
        when x"FF4" => cos_16 <= x"7FF9" ;
        when x"FF5" => cos_16 <= x"7FFA" ;
        when x"FF6" => cos_16 <= x"7FFB" ;
        when x"FF7" => cos_16 <= x"7FFC" ;
        when x"FF8" => cos_16 <= x"7FFD" ;
        when x"FF9" => cos_16 <= x"7FFD" ;
        when x"FFA" => cos_16 <= x"7FFE" ;
        when x"FFB" => cos_16 <= x"7FFE" ;
        when x"FFC" => cos_16 <= x"7FFE" ;
        when x"FFD" => cos_16 <= x"7FFF" ;
        when x"FFE" => cos_16 <= x"7FFF" ;
        --when x"FFF" => cos_16 <= x"7FFF" ;
        when others  => cos_16 <= x"7FFF" ; 
       end case;

   end if ;
end process;
end Behavioral;
